%PDF-1.7
%����
10 0 obj
<<
/Filter /FlateDecode
/Length 23
>>
stream
H�:��� �����pn@� 3
endstream
endobj
11 0 obj
<<
/Filter /FlateDecode
/Length 2818
/Subtype /CIDFontType0C
>>
stream
H�|TyPY���+fh������JTtaF]AG�@���G9�
����@ @ 9"�C� � �*�
�Q�x �%�:�ʪ�[N�v�-���g��j�������������ǁ�@gy�����u��D&��և�SU��rGq��+*\	z%��hM������
���ޯ��K�h�i?W�KĮ�U���z�q��ɒ��Db�R���ek��4%�����ˁ���ى[��͉�^�fooo'nv�ʩEEhJq���'M�ɳe�D�X����̤��
J.V�幎��ġ$
J,Q���T"[L���r��R�E�Dy%sT����+J"�X-*J*q�%����������,SI�r�X�a�ވHM���D��.;(-���\h-@�(��CP�p��!(��ul��e�2�dàph���wY��w3��E+�xB>���� V�3�Ղ��Km���9,z\���e�B��
�i�w��dj����G��P�p�N�8�`��,
M�1��w����O�;s�E�:/]ſ��m��5R^us��G�\�)e���/��'u��!u5�r�ᘾ���������X��\T��S ����'�ȓ02������,hmm8݃=�����L�p�'��s`���ʺ���� �oᯐyZ ~C�ךf��pja�Lh؅3u|dF�����x����@�@<s���
9�7p����c���&��Ҁ�����l"Lu֪Ny1>$p��ƅ�OGG��<�t�cu@�_9y �u���B;���~å{�5�Q��8�Ÿ�� x=��g �qt���1�.�/��Z?��ÐL
�	�0��ɩ�m5�dK_���4V���s�<��^r��c��ӆگ�b���Α%����U��}rzb�)pŞ�ݍ%&���g\<��������V=�ߚ�J/����7{`̖�ń��> ��+�e�}4�;G;�� ������y�|� G%���M;ѐGj,��o06��ư�B��H)?��L�	_��ޓ'��S]��FҢ�S�{�?2^)�݉-��~�P_k܄-|��y�	$WF���3m�M}lpCa?��?;�J����(S���c�08Q�U�%�L�g�|�v���"�Y?� �v��&�Ͳ����5;��8�bxL!�0+A��#k������l?6OVU�0�4��n�38�Ms���R�PZT���5M�Hp+���C����Yxx�~�L-�+*.)Ĕ6uKc}MsQ{�l�XuM�m��sI�I��d���y9�q��?���wt��Q�o*�	J�ۏ5�G�4i�9����1��u��l�mo�c����Q��Y.�.z�p��(�5ȷWo���zI���X��[���Fsq=i)H�$㢐��h2(:=h'F���'�	���{+ao��h�D��j�󿂢�N7^A3*y)U��1�~�F�
x��ڸCژU0b�UJ+�pf#d8�_L��m�2�$����Èl����Z%@���IT�H-H�L�%�������i�0�My�pf@�.��*I$��V��`I���T������{t�7:*�p�tD~h/��� �3wZf~ �`�z���r��`���"�#🛆�Fp�������?�z���֕@e�y�j����'[���G���_):�ޏ"o�TC�!� y��,M7K��?���Ky$��h�:#'����2�\h��T�K��Q�Z-(,<����O|�pq�,~���_[0��>��Z��Ѵ�56�4����-�S��/c ���ɳ�׍<����f37;��%������E��r2B|�����aҺ��~C=��N�G{J.������.���u��	�g�XM���I���;�o��>�z���t�c���UYe�
UVv���F��P|��7���K8A_�c��Fi�W���D,��*B��j�73 ~��ۖ��0SY�����]�����<_U�.��	�x��Jx��d<�1�𾲲@=��lp����"�@�z;/�:��%���z]��Ѯ��>��3P���t��,���1�G�-����4�7 �1�5�.���j�,�	�X]M9T������$�����?׎w����I����[v_Z�uă��I�cI��M�q�z�>������Ká������|�ȑ�����������s�i[`SYm ��!������������ƃ��vp�b/OPE>�j�o�t�s_aiofO^��yq�g�G�}|��x�����X�@�^�c��������cP��=������������}t�rrj�������������}�JIB]pn�����<�cʔ������v�;���0�\��q�I�FrĄ��|[uJk0h8n�c�q�{�������ar�����Q���������)���֦ǔ����������!��6��A�5�!��o�N��f�)�(������ԯ���Ȓ��Jr����ykyjwlwnP�y�������\r���Z��n^pcoh�cY��M�q�O�W�������������	�p��`�q|��v�1���3�V��r�I�Iră��evL`�
oG0��~�������_r�~�T�D�����z�~�|�~�vxht_wrlwz���{s�s������������4��9�ޤ��Ĕ��� 
�&�s|��I����%���������F�_	��
��w�n �U-
endstream
endobj
12 0 obj
<<
/Filter /FlateDecode
/Length 304
>>
stream
H�\��j�0���s�{�Dݨ-�P�]�?��h2n5�����3��>Ι=�O�sc���&٢�A�p�nN"�xՆ�(-�F�-��2��e�86f�XU�����'5��g��)t�\aw9�{�����xH��A��^;�֍<�t�C��s|-!�����I�l;��3WdUN�9���Q�����~�ߝ��4ؓ$K�R�x��#���4�i9� *��H��99r
r��L�)O��Dt{I��YRfN�%e�%QA�H���t�"l�=˛s�����ڪ6x߼�,���a� gɘH
endstream
endobj
17 0 obj
<<
/Filter /FlateDecode
/Length 22529
/Length1 49584
/Type /Stream
>>
stream
x��	|U��7<�9�InB��%���-$!숒�$� aYH0[��	�	�

�I�R���"E��E����Z��B��H�"����~gν�M��}�������;s������onB.���  �8��3�W�v�!��Co���I��߫(#da��9"#�y��O�����Q	��YB��c@pocW�.�G}�G�g�M\7\�*"�?�3��ym��NHǋ����������Wq��잚Z&�P<ۧ��_��{%!]B�%�e�\�i$��.@���a<��s���ʙ)�T�xl=��4'{��K'2x�s��g��0}��K1�Y�]������ލ���J+*]�xBԈ�e�ye��8��jBLm�����s�-��7�;b&�z�x��=���Q�������<S��:���rW�zDb���ӝ�.�q�M�:t%�]CT��P7�1ظ��I>��f�f�1�o$�����A'1qd~R.�#N�K��fS1�|2�W\W$���}��)4ԏ���s�]t�I��Z�K��|���"�2�V���,"��5��d�r��!��#N1~9C��'��[��*�\A��Z"t��[��$��#�m	�������#I�,'��YF��K�{�����?��@}p�w+ț$=oЁ��Kf����Ӯh%�d�!fO�+���5p-�kॡ�9�.g��,e��x^�.�x{�7��n)D��.ˤ��-�p�HV ,���
�z�e�cF=u��ߤ
:�$��}M��媅.bL�ih�����zS�l' ��:���հ�j��R�5��T1�nU\�R�-���� ǁ�װ
 � 2����d���ed F�$mI��G����R#N����\-��I���c!�P���C�-(�Q��ß��8��8�Gv0.�/�%(ލ���V"����z	le��R�b��=s��v�mϼe�@j�Cţ͹d���Z��'�C�����B���4�8�gJ�E��Xɗ0���c�5'O@��c�s��Gg��P�����4>�ç�w>A^�,�nCL)@�
���5��DvnDɧ���6��0�e:,�:��!~����sxS��Q&�����b�~G�do;��ވ�������!l�tO�x�/�&�it�Ok��(7���(�igց�/*��r E�{�.�ь��t�Y�oh8��i �Dz
y���-��B�G�3��h���t4y�F�\�� �%�-�����������-r@�[E7"��/��[�39WbƕEVF3f��#V >���!�X��U5"m1�$��5W���+��G����-������#��H�-cq���3�V����Π�����hm��Y��M"֠��$�UI��w$֓�@[12���=��er�z�
��H(�a?�NAmy���1��X�
�n;�<� o��(�W��u���X�Ů�I(z�)�N)_{����B.8<҉=��$@��x.G�p��N�8��3�\�>��OH�R��_�uBr�)��`���K0�Ÿ4�\%a�ki�ܓ��'�('F>�ǘQ�K��@IhTĆ2��
XE<��p2A� �[��3��5���7�c�ϖՃ��ߊ&z�䩡���x�~A��2���ߘO��i-b�C�[�,h�Q�P'�g20L���C�k��8���ce�Gg�O�,��0���$6��6�	���%���U�;��J
�
_%�`���W
0���߸���Ndua��2��=�!��t%�U��ڊ��>FMrg!_�/]�P:�8\X�*"���u v0�Ad!���o�u��Ub�eV�z�b	,r�GQ��Ӵ7�?�I^Š�%i���z�HvS�{~5y��Yȡ�lR�>+N#�d��A�Cq�M.ޗ�ga�Q��������u�aĺ�$�u���B�h���m#�bG�#�Ϻ�n�m�bw�#����b���7��V���[+��a���m4�>�{v��=��K�֒�h�T�H�V���D��(Q�z���xr}I��t0Jw�(�i
��;3�P��g8O\��Ci��0��X����c����x7�f�`PEĤ�bV�l���әt89O����1r"p� .��Dvᩞ��S��ޙ�5��dT��,�kv�{���ƹt[\_�fsF�:"��M�z��?�M�-��O�'3�;/[DyA�<K��R�ӓWx�wn"2+�*h�|ʻ�Q��d�z�^�j�2�^s��������խ�[���n������^���n����`��F~��H�a�sw��s�=���z����rD�FE��IzPS>1'_�yY���o�K�{��/����{�]/�ge�Y~�F�]�#b���`�����
��x�kp't�����W��~�u��tV��#(�.��b���������N�[d(2����p���Gq��Y�Z���u���:��1f7mA��8�������c�8�*���'yRB혗��}��me� %=����a�#u�Ⱦ��ḋ�1Q��h�TWhD�.�����8�^L�;�Lu��ޟd���pv'�<��cs�����ڶ�V�K�X��w�mϓ��
��Q"�>��^���-ka��}0�]�.��o��>�.�o�މ�V�[�o���}��-��(Ȝ(�u�u�,@Y膷�`��7��]�	��r{
�<��w����g���K�,hx�gg��2�Q{(J��Iw��.c��i(YM��,�P<�(#�(#ݥ�̶rn!��� ����{�4��|d�A��<R�ROy�X+��p�#*Ff�O5��N2�dA�mEeYF���g4���(�����i�zzý�6z20H��h��O�v=��tS�ވ5�ho�}��y��i����F�di�n�V�v��N����l������jX=��~���	HO��Ƙ�?{���U��᪡3q�Igz�޽}gaAn��,����
$^w���
�x�Q�œ�ɧv��!��.2�}�����X5�'z�˜����Mg��<��h�§CA�!>�'�Q��\��>
���s���-No}�#PE�ELՎ��i8���s���3X�`D���9���I��X]{pzHEv�X�����sx鋷ca���l�󦁛u�3���ӕ/0��dhý;�����h���d���Sw��!S��.
|E!�*Q�g��8�,���i��8���\�[p"F��=�*�'a�n����g#f,�In2�8��{�38���}0��Zm	݆�$65�~�(�6c:�},ƵF+r���h�@	�'z[���-�SD����ҕ��o"��}Q���B��B����ͧ%���;(o����V8f�JY�!.f ��g���ޛ��# �9��:{���$␘U�w�ω�f!O�9�hgډ.�KDf��"��4hv�*�FB��)�1�#�# ��⩫a���?M�R�g��*>?ނ�G�'��$��%�f�N� �)!G>�K��h��͆���s�&vk����u�5��.O�?q�w����Z$�=�ޮKF�qG�V�9r�'��CET�<�Ơ�F�xB_�W��q� k晇��Z����;��1>�4��OW�ɑ���Oyߑ�6��&���z	q}-�f�o�}$��d�G~��y�,y\�]q$��	��$��D=W:r���&��OJ����I���,�ۈO'�Y�V�����g�nn���5��A�i�%����I� �C���L���q*��	W���	��I}�T�sw�I�-0�8
�#��:�"��BR�h;�v���\-FuBD��Q�UB�1��\���w|z����~�%������s���Q�|��*�?��jC��ꐧB�g��P�&�F�wW�>�]{�I�Q�C���*��55U����E�:���A�r�Y�����F�NA~��⇆��`�[R�[w�������~��ܭ�es�Mh�_������ xJk�m���KN�Y��:I6\1^������w�[�F���ˆ`��}5U�:y+O�v��D0+v������3����px��&MU8r�H�c/O���`������"�<:&�^2r��,g��52Ki��ݫ�����{��O���"���rVӖI�n�I�љ���xB7���;Au��)��:s
�����/w����
�O��[��ߖ6������f Pr�/�	��f@_������j|8�A���!�SN��E�2#q��$ۚ�ʶ"���a��ƍչ�󺹼V�?��v,��!��\��[+���_ǔ[ߍUo���+�݌P�˿�SnF�o��V��Ϳ�������#�_�_��5`�F�5ծq.���W�rկ��k��K���6��t�E�W�_}�����O?i�~z�Ҋ_Y�?��_t�ч�Տt�as~y=����?���U6����������.��u��;V�]��c�t~^�o/�W�n��j�������O+��?�������u���_����>�I����q����c�w,���#�R���������W
W?��)���A����W��W_�������:)������{��:ߣ�����|���w����}�b�������s��N�?;���3�������:��ηmm�n��[�u�[[�g��V�E�π�3:���7m�R7�|c� ����OR���i��Ӈ���uk��u�uq�Z�?��'���!�&���2V��' ��|���D��\�J[Η��e:_���u�d���D���c:_���	���@��g�y��U���ѹ|n0���G|�l����t�WU��*?^UMI�e���+�)�"N)���t^��Ғ�t=/)d��N�H���i:/�����C<_�y:��yΔ`5G�S�C�̳u>Y�t>q�M�����N��x���8<:+����h��j�J�3u���t�?8�����@���ᴛ:\穇��N|hJ�:�O���!IA�����\����C<)�'�#���
���Y\�EI��S�yB5#x���U��x|5=����v5Η�U��xh���|`5���U���`���|��������/����Z�;���y�n�jo���{ƴV{�=p��X��yw��ޚǴ��hE�(K5���L�ȻU3A6��F6㑂��J�.�jW�w��.�3�v�y'�w�y�o���'�~<L�~~j���;����rg72��r����-t�V�m`�6�xk���y��[C�dޢy7�Eo�P�w���� �й?$�O�Pp�s��;?_��������XU_;�5t���X�t�_�[�]�VŦs+$���҂�ܤs�5����C8~�C7����n�88����WѮ��\����W;B��鋺�>�{>=��y��<E�6��p���2z흤p��Z�8,�)9����q3W�*~���3ʇh����K�%��`[�@���ߟ |��Y8a�t0>��dÝ���7�p�e-�AJ��-�!�qN�I6�k����s
���~%z	Y�<�����������.�ɧB!��u�z�u�����)d�zI�(��%���N��Ma�B�m'=L��4�.?5������t������jF�d���V/i�d�)�����,e�,���e2�E���=���������ijdΗ��$�jj�&��?�t:DI���E|~�3;B3���^�^JQW��B馮��_j��`8��|��ނ6Ky"����d1���i.�Pqf�|��^)Pw _7���2�"8�fu�o�'/�t'��5kb����o�߾@!��M�_��&��)�d��h:�š[��B8]���f�0MQ�@��ts@Ml�����sa�z�v�P�K��Wić���i[�3�>&�4d����~����&�j�y`@˰֫g@^�xѢ��6�[�A�����_��_\�'>�BO� �����kxM�f&AJ�xkkb��h�<���z�����s�k5��+��j���~����ͥWx1[���mL�Dq\<)5C�7oOs���_l���%��.��d;���X�$Z���jkiw�m"NO�]�+��QNHa�ך��%`C�}C���M���ړ6�~��C:�iX�qD�����������8�G�h%Z�֢M��hK�5�6���@>P����ZZ�F�taa�D&�Il�u�m+�J���|��Uݪm5m5o�l�n��H^�/���ʋ�ڋ��/Z^��h;J�ң�(?�U�jGMG�G-G�Gm�?ƌ���LR'i�L�̓,���!��}����#�E�@-,4�Y(�w��w��������}G���w��U+V�zbŊ'���w���͛�z��#��MKe[�����~���޴�٦�����t)}�Γ�)L���������@�Aaԥ&��bӂ9,c�O�J#���D���_�ޗ���Бgi��ӻ���꡷/�"�F��}ے�:��᪦�j�[�	�45����φ��
����ʨ5�e��wh��c����	�<�#�ɡ~�߲����ڽz�>�^=#�B5S�h�X:3�RZ���V�A�r����l��R��ܾ�v��u�F=0{È�O$:�=�ګ��UƋ_�&���}�o'2�6��ܺ²�g��¹�톰�ڦ�/tnь��V��`h	�~���0ﬁ{
�u�q�_��X�c�`���v���F#��y����M}oj��Sv�۷q��[�\2�H��WS.Su����o�=�Ù^=ׯZ�i���G:u:�t~��Gv��$�B�vd� 	q!ԇ��}��6��/�P��������Q[{q��	P�U�
�g�Y9%�j��y��Ekߋ]�;�����g�W�����Y�c�����[�u�v���P�Ԯ���
��|���g�iW0&-��5�8B���O���U�������/�B��F��z�ݬ;�uL�ԡ����&�~�{p3�w����O��U�~��|3��������C�8D:��0SH�֐��l!O(Z�wl
&>�&�-m.�M��#ڀ��:`Nسy�O0(h�K���mAC��-F���O?�z̮������F�����`ݺK�.U��_�������o��o�*�$�MW��ܱ��~�g�\?+`�>ЩFzŵR�g<\Q��*��4�����Iأo�x��cC�K�n�����]f��^}{��U��E�I���a$�������6 �v|!&�ޡKp��~���mBy�_����F�Mh����t㥂�(,Kw3��@�4��1Y��k�^�t����O~s��7O.X�Uׯ^�][�ϟ5{��Gf�g�6,_�i��e3��}���oz�٫���v�N���3g�_`��<Ȕ,e�@�m��-~��Ya±!T��v}��f�!��`{D+a�5��gS�~'��a�p�����؄{8��C#X悵ka��?�>-����T�F�����ul�ǔu�`nڞ��}�Zo��Z��z���^"�	�_*e>�&·m'���J�)�V��7���߽���*�z?���Z�S�p��B�㚙�k��d����Ҏ��iV��(焠�ؚ�f\�U{js�v���tC� |/��Rf)3�{��T�Q��=��M��NJG�t���7kZ�����Uf����?\Q����c������t��K������2ڕm�F�*5D<[�{�����\���
��f	��� �v�m[���֭^"�Zl�>/��96X��M����Iw-���a�¢1ᰜ����{����w������O�t m7~��F�:y�T�)�:w��i-��:w~��8l�o�o����~��2��L�I�����R��O#~��w7;b�H�����w��wD��o&��L��~�:{�E&���4Q?���/�����~�a�����c�~Z��6�z����B{4����T�t7!���ٱ	zR�z}�z�O��dOԕ���3D�L�U��{��*Y�m!⚹q+��$�V�!�7ڰk��n˫{�O�]u}$���7��dq\�a˄��2ja�&XM�3'�m�Ō3�j�4%ڪ�Cib���D�����gg��g�䡸��jiI�xKs�%�v��Ζ�8��6�����P��T���ʰ|��F#ca�~��[���"37��owU;�~͛����׆��:������3_[xpH���L����-8D��_
|.h�?}�<�l_￩S����D"����h��I��ښ��e�#4�e�h�FR#o��(}(�j"&
5�}�<dl:"��%���"�v@��7'�2q��⧧�sL������ol�U�d�������#��7���W9aA����O�u{?%q�#eӝ���l;�ώ�= �;"����a�p��j7�m�f1#�3��MnC,�2U�8�'Ė`3�L�i-��lR�J���hr�5�y��j�i�������M���>L����؂Ԏ��Fزl3�,u��&��~f?s kmn��ծ�p[/6��5g��Xs���P��?:��X]i���?�O�U��M��M֣.��[T7�����J��.'Aq6��@�	抌R"蝌�h88R��z����Z�3!��rA/�<�?�j�7}�}JB��\�!Z/9�ثDN��4�3)����vڃ�L�@�ie@�Σ�Vv8�)ȇ)�|��=ѩh�肐��5�r�'�ެ��ޏ����ĵ�	�qƴ�	�F��ml�u�m{�m-�mk����Cng!�W��^bk���|�%��J[ WcG���ogm�C_y得�������.Y;����CY+N��d=~U�W���Ωuv�Nzm������ݳ�c���ص���A�,��m8	�ĵ�[�J?������y�	d״��� [l�qА��H+<;1��2�G����K{��K/Y�|��u�G>���k��U]͢߻�᥋]f3ӳp���w�Ԙ�U�JN��p���km_�s�AV�:�b%w���I��hɭag�^��o���.��G�J��_����4�*nNKY����=yc|��]i_�ҷK�k��?9����= ��� KC/*	l��7p�y���o����z&o��H��Y�[�q��Q�r�t�y�u����X�x�R~��wͪ�1�>�P�1���]���e?Y�Ks�AZp��*��������Z��Ϧv��uXZh$�m����I�U]��y�(���n�4�h4n�d�~~tOֱ�������y�U+O.]���&��^>ݷ��P^?ڌ�i����/��"��zkFzBkj7��J�v�ʚ��E�|�l�"��Ez!��X����#��vT�`8ش����B�p�@�W�_�]_xI���Ԝյ�����=�?�Q�kvH\�V��6-<`E����-V�q��`���w�؊h��Z@@�!X�'���Q礱X���5��f��!��ϼ�۲W>���?�z�ǫ��-ugƔm��^����W_�,Z]������o�����_j�ڶmDEn�k�;q�OM�L��������������r�ӿ��G��`���PD��@��R�-����@�`V��2H(m^���+���?_�؁�����'^�]��Z`ݎ�9�
���Dг�\��|��OZ�!�5v@�6���d����!`|��NTe��)k%�}Z\[B��OiHu�2�6z�j��]rm�*q�,�[�O�*װ�l���Z�9#!��Y��}�"z	?`�Ə}����Q�3�B��yt�����k<��ݛ�����u���j�3�R&?/�%�K��!��Z�0dd+�J��,~�<��Ar�y�-�N^����k֬\�fͪk���յ[�����]���K�]ޢ�����]ڍ��"J�=��V2AWģqm����M�?��h��J^�>]����t��F�{�+�����/��o�77�����h��c�����ό�߹C��U:�_���h�d�ğo�=b9nB�H���'�	L\<'����pqP���8��?����#qt�#�$IG:F�<D���`��ʢ�f��> >�.J�ޛϊ�����w��Θ��X;�`�t$Uqq27l�N["GLh$���d=��h~,h���2���vFz8���b�C�:��Qz�п;M@K��{����i2�y'���s��o�ؖ1��	/]��杌ӦΜ��;s�֧.��S�?*���aC�|[o���PXؑ^�r����|C���͋���{��,��{\��j���?=n>`5�,���mekn8)?f����h}��|�]�8���O��%¬��~|uݶ9S������>�ޛ�(���MVz�.��P,8��j�Ǻ�Z3$c	�o�'�.[���W��������bK���a��ٹ��̅���d�s��:c�EB���k[r&~�����q$�ⴢ��$�<�J�wMd��v����H��ܬ(*g̓�Ұܣ4�&�˿F���f�N�r�ة\��&��*NN6+ز�'��	i5�4�M�?;��$��ʸ�k��l�Y-f�7]l&}�ȸaω㎔g*��z��V�,�-���v�5o��R�Z�X[�B�'-�v�:��̑�~���O�g�a`O2�X�mC��Y�1���|V��Bu�%�6��Vg��X�m����X�k��+�>�PX�X�Z��B�����g)����<k��ߣ�h���8����O�o�}i�^(pK�;�����m6�
].�.m䅸!jKͤ)-�b7U����Y��#�--V*n6+�ki	�〉P��3w����$;�k�I�!��/?Ę�F�-T3��B�t:ˤ�|gҬͭ����q�h�2ZX�<��E��z)���W�\��z�9ڙvT&�}YWM_��!,H�>m�Z��� ��mqI>-}}��ؘ�����2�8Z�9���;||}�Z���$8��_�J�	����~>��`H�Mj&���r������Y��7@�][+��f�7����������0��*β���|��!x!)��9�Q�'�+~p�`}�	�J��UG�����m�xRI�]ǋYe.Y-$4. ��;�0r��q�jM�O*������5Ƚ6L|Ɗ܄�4��%�҂���+v�<�<c=�k�,�B��D�6Kj���XD>d�F�=��]$w2��'>d���5E�)~ث���|^u���9���j=��������3����W�I��kN��� �k=`�Hv���Tin1!HYl&�!~I�>I-$[��z��������^d����/���Q3��8��/C�J���� ��9��f����Cܞ���J�R�lV�)�5��:E]�V{-ȫ��S����e(�1�ٜj^g������r�rS�%˺����c[�m��=��=�~ۧ��{��{׽��u�wݻ�]��{׽��u�wݻ�]��{׽��u�w��xM��~��+��,��Է�orL"���A�OF��������~ū�;�p�5�K��ⷵW��6Ҏ<�n�X֒w�m_���Pł�#�<w��-��f�l�ns�~ū�� �0w[#mm9����6���wۧY���n���o���*/�ZP������9e�3�����</�8ҙR��/*r��Q�������y�Q�ļi٣��9�%S�*���y��gYՔ��gniqva�gLFvI�sxiIiBi�ã��+
KK��Q=���k��=:���*A�����tt.��WEU�V���嗖O͋*ɫ��Q�pataIn�̨���������d9[p#$���٩"/�9%��tF�(�/�=�jm�����z�Y���e����u6�\���ٹy���;K�b�ZG�VH�btA^yhM-�.��ˍt�CxL���^���ԙ]2�YS`B�J\X2Tr��YY��6DvNNiq����^dh��)T�$�3��:�+*Js
�A̩*�+�̮��AǝF9��Q�_9:�,9)�++/ͭ�ɓhr!Xᔪ�<�C�	��RNQU��dFaeAiU%�).t��UmU�q"��yRjiߊ�H/��fti��"v��B���	i�Ж	EW�U'	�((-�s�0C~Uy	�ɉ��Ί�HgEՔiy9����q\R�SZ�[(��o�f�U����yRË$�NPRZ	3T��*e`�sVdC�)yn��8yv#9KK�����򼻊�U���BQS��g���Ks���eU��� ���\)��:�����WUQv�$��WQ8�D�1�hVYA��$<4;H*�?M)�k(,��A$�y^0�Œ�Y��F�����7�ȱ�Q!�)l�Y"y�<C�������*h{^8C���j�u��	�`5	�U��bzia=cy3+�j��eeXb�S���C~`nb���JgAv0�4��5xx��
!��+�q\	5$�)�V���-M'��,��3�,;���k���>~�r�jD
A,����$9�G�e:3F$g��OOr�d8G����������sh�sLJ��2����9�9"��6�9,%-1ҙ�52=)#�9"ݙ2|djJ�R���JLI�L�����Ԕ�)�@�9BNu�JI�Ȇ'������Ԕ̱����4�3H�#��3S�J�Ow��>rDFp$mZJZr:�$O�@4h�ȱ�)��dFbR&:#����I��ӇE
G@�t�.�Ù4ZL����LH���LO�.�
�N1\�hTZb|fʈ4gBD�OHM2x�(�R�S�G:��N�h "���iP��08)-)=>5ҙ12iP�h@�)�I�2�H��H�������(t`��2$I�� ��7Hr&�O��O���zVƤd$E:��S2��#���'fGA��xin~��DߝށQb�[�Ĥ�T �l�1ޕ43'��R��{q�Q�R#~FJ�5� \xp	��'��g�,���aq�-9�~E��wc72�o��<D�
J�>JE0�QX!W:���R��W�]b�U?
�2��*��l��<bYy!��(/�D0qfW���p�{+.woUM%T��_�WQ���pz^Ѭ(�-��䤰YX�[t������Z�*��Bp�jQN+�d���"夐L%��8I'�C:�KbPz�5#�$c*�XWbt�&�$�)���ב�8Iz=�
���{�L��H+IDk0�&U�����2U�t�-�;���c� o!�91�t�廦x2$�a8F��&�����^Я��R�3\� }�����m�;_�U��V����O���O��(�+Ž\~兘[.���<̉&3��è�R1w&ޖg�R��y��<��Eۣ��xW!�@��[4W
j������=J�y��Q6����7�w��U�������;���32���ﳥU��VF_)���x�����%��5p�wyn��J*%�s%�|�6���aa��"%_���9�̽*
��X*�.�^aȒ�ִg���Ȗ_�"<�̍݃A�6x/j���Z�^^*-�-ׂS~yL��#ׅh�>��,�X*��~��K5��S=�Dt�Wb-~.(6�D����J�䳁�\)A���)x[)�zh�8�H�Z�gU����
d��tk�X�yK��_��+n��#��#��Ҟ[7��
̎�9"�化Q�)1���]��jc�����ܖ�{te�k�h��G�/��Y�2�%��+��)�B�0"G�3�x�q�;Jz,�#i�J�ݜ���3�=+Kedh��w,j����@�.���P�h�g���5x�sJ��ݖ�R�=�fhÈ��?a�R�#9ݶ/������b�,�o��wT#M��\��Y����W(ײ'�	�+�Q��18:������y�/A��W�d�y�r%��^%^ژ*��J����<14[z��M�S�2yǸ�F�-mt7~�������n<F��^$��DT/wG�<�_q#����z������H�;��5��)U��z�}1�^�3�xϮ��m��Im��L��ԋ�*�z�Xb:��Ec"'�t�5bt���e�ȚW?����?�b
d�w�{���<�Q?�/�tw���m�;���W�O�+��l�߮�
=={vê�(�A�� ���1�I�~p��bƾX"u�4���"b��TS�k�ҽ/��kjI�tF�4<	:#�I� �L����78�ϥ��h<�?՝(�/߈��r5�A[`AFI\�t@�{,zn�|O�0>���$���b��:m�{8zSqOr�3ė{�³h&"5�aV�\;b����4�Ts�")z8��t��~/�1U�+�'�vZ=��nN㥎f�s8J�O�w�#1.C�3^�lp�&eH�{C�$Ɂa	��A����ϣgJ.�L��H)��'Q�T��^��n+�v�(�.>��G�Sΐ�8����ɔ��~^�������()_���I!A�Z�L���e�AR_�n��DI)^j$㮒x�5��ݼ�Ca��/Ij*U�΀�0>�����)� �n���>���ARFa�A5��S�Rw��0V��A
��n8�Kg�Os[wP��GH/�S+c�ZL��⥭3교,��p7磼<�c�Qn�Q�Yc�z֑g�/�.��L�����0�^?�׈]I��r�y���D�k�s{g�Y�w�Ib�w&`D��rlq�q�F|6���3�ww���sJ6r���ד}��8yg��2O7r������?J�3��mÞn�����^��kHV����_f�lAP���6j�jzB,���Ae�lW�3!_�{����T\��T�s6���s�/��.#ƙ�PjX�Qn���s>kЉЀ�YXq�7x��֟4�C��zq�붸񹚠i5~@^�G�w���{N1�]*Ʒ���>��oE8{�P��mBk3ی�3�7hog�E{{��.��^D{/ۋ��+hd��~������O��h�Q!T��<N��Ty���y�/(����	ڟ�>%T~��]��H�}��e���>1�R!�w�~�d/��h�ɩ�$"�<{
�əU^D�Z��0Y�]�$��+Kp�U�&\�7#������ �>�д���Y�$攌�N�s����
�&��3}�3cX�����*~J�FJس���I���)��K�����P#&)��K^J,�	&���k�o�A�Hw�g��6��f��2�x�>kh1�6��n��;XR�}����(2��eeuW�le���L�c��"��`��sX�)T@��-2�Be1�\���WI��&��tk�zH�V�H�����d&��/.��U��?�����OO���n�G?1f�k)ƌt=V��<�κ�Y������fw�@����}�H	U@GM%�Z�c����UC/�O���~C��:S��9X֖��N,��d�YKf�,�e��,�Mcel:��b}>��a}nc;�n��U�#�$;�γ��G�3�%��n�ۜp��y �����cxo>�'�!<�g�q|2��E�������r����[�v�<�������������*����x����*���D*�J_�%Q��TF+�)J�R�T*�a�%�J�)e��C٥�U(����i�-�rY�D�B�Q�Q�WtUQ��Cm��UC�Nj��S�Ʃ�j���f��\u�Z�NW�ե��:u��Mݩ�V������zV=���~�~�~�^Wo��5�i�]Ђ�`���E��zk�m���ej��Z�V��k3�G�Ǵ��m��Eۮ=����k�c���9���c���vC��՚��l�5�Z���S�)����)�4�4�4�4�Βϭ���戶k��]xa��3V���@Z[wN�V�y�u/�]s$\)��}"a�Đ
�M^�I�Щ#��LW`�k&ޮ�ؖJl�e� W"`'=Q�r��ϩ�!U<�uu+�OY��_@I׋Oֳ�K�ӫ?Wre���|+�fI8D��у��}.� y���=S�ɮI�>:8g�u�&K8��r=\,{�$̔=J�%{�K� {&K�PbN�p���q�-�-zR$#{2%4F��p��yH@p=�u�8����h�'���K%4��HX)9�  ݭ�H�%a��"�s�ș%��߷�9�WK-�d����޼;d%W�K� !tK�ߥ?�i�l;$LV��-F�ۅ�$<�A���9	�\�?K�K��k����&�+%�F
M�"D^��
�|LjcN}��y���tU��5��,׎]/j�O%�����h����Bz�N���u�ַ���z��Ro�H���ڠ=��߀3�@AK�oҟ*18��+�~��>/��oԷ?��f׽_?q��]���?��*��MZ��Ϻ�О�Z ���{���`����a��zPr%v����ѯ����r<�� �s�.r�dWsiǎr�(��u�Ě��S]��X��X��{�H�{G�����] �ҟ�S�{!��믯�t�l��fF�I~Hoʞ�2�$�H���`"�0⣌Q� �/3��s$�e�a���R{'{WRa��~�aO�"3���]d�}72�+>�>��>�}:�k>]}"�W��N��e���\f�&,��ԫI�xS�&=Ϙn5�)������M�\Q���L�=[eOC.cA�>Wfl�E�c�b��ⷀŷ�ot�E�� 1��p(��c��I��N8厞���H�S��3�:=GߡЏ�U��Ao�ZƘ���@֚9Y�d��/{�%��l$�&�)����J6��gK�J��Ȟ�YeN'�av琷�Ev�}¾`5��=ӹ­��[�<�w�Q�'���x2O��<�O�|/�����/�O�u|3��w��|��G�I~������g�K~����h�]	P��`���E�Qz+�e���d*��J�R��+3�E�)˕5�ze��]y^٣�W*ǔוs�;����U�+�rK�U�jV}�@���T#�H5V�>�&�CՑ�hu�:E-PK�Ju�:_]��T�R7�Ϫ;�]�^��zX=��V�R/���O�/���{U�ͪ9�Z[-T�Ei=��Z����j�Z�6Q�զie�tm��P[�=���6k۴��nm�V��Njg���{�G�gڗ�u�v�DL�I�J�s�"��W�X��jaoM�n�VD`e�~��hӛ����"�#E���؅��"sP�,�Q66��@�#�if�S�x�6��.�H�v��zSD'%�V\mQ�G�9_���܊��+"���Y%�g�2@��	�V�]� ��# �$��[������(Y�1^p��qfz����0A��.�T	ǫ� ǩ����0EyQ`�=��*��(�0U����Q�,}��B�Z��d�S�¬\��"����A	wKN�d{��;%|����o"���]���l�g��p�C��.���?۫���*v%���O	W
�o%����@����@Z-��>�# ױG�3�K�{����"o�2��b�:R��G����G�r�!�����|�]�?R
��m;?-}o��R��#0�(�"��I������j�����	�/
o����'�)⛃N��Hc�5��Ǥ��,�Ud,N��)b��+�%'BF��$��o"��E�N��,�~"򁷸8_����-?%�� �U����ugW�|���� =�7�<��$p��8�t+�\T*E�"�F�iɕ��l_���/�7�V�i�� }LR?/0Гj�����i1R^����d���}/z���X��U!u��A�U�a�rQ�E��,l�fَ&�~���ǪJ�
���bi�2.����k��"J��0��D�
���y������j:z��`�|6�/�hp��ly�~Z1��d"���--c��ә�l�Kx/���������9�Xer�	�d���7$'��H��t��L��g
d>Sd�O���d~�L&��ŧ#�e>sE�3�����-�Xc�.�Nm,����a�� ����4��Ʊ�,��r6�=�c����ma���l�/>gd��s����]e_�������@ޚ;y�䱼/�'�|$�'�)����J>���K�J��ȟ�;�.�����q~���/��������﹮(�Uq(-��J��I�Rz*��8%YIUҕ,e���LSʔ���Be��N٬lSv*��}J�rD9��U�+�))�)_*ו��m���jW� 5X�vQc��� 5A�����8u������L�Q�1u��F]�nQ��ϫ{���A����zN}G�@�X��~��Po���̚���֜Z���j}��Dm�6R�MЦhZ�V����kK���S�F�Ym��K۫�kǵ��[�E�����V�}�}��&�d59L-LmM��N�(SOSS�)ٔjJ7e�&�rM�Le��������0�3m6m3�4�6�3U���N�ΚΛ�3}d������鶙�5��`2�;���c̽��	�!�43����M�$ �)۳e{�l�?pJ�g^#e�{��n+�\mC�4�Q��w�1(���sޫ=������x�}E��ƥ,J���Z�:. ��b�o�[Eo�,o�~:��=��Mu��Ҟ^8_�y����'�xk���Sj�z����K^��O�{7է�=�K�_����]?�6|�=x��cmH����^3i��7'^m�_S�	?n��i��K佚�\Y�)4����=�[{?�����#~�����^=F��|����s�xe����$�����!K�z�A'�4���ľ���o1����?Er5����qGD��iM��IO��l$��f�I!�H5C��$��$�H)9��+r���������W����|K�&�ȿ�r�ԒM�E5��Zh3����-ɋ�5!��4��L#h�
�M&o��oH�I�#.v�]�����9�l/�^�ܶ׶�*��l��j�h�DM��mW��_֔�X���9B��Ж�	����_�3�S���Ti�m�oZbZizʴ���i�i�i������-�E�e�'�/L5�oLߛt�b�����Ps's�����9ΜlN5����͹�i�2�t��B�RB�O��3o6o3�4�6�3W���O�Ϛϛ�3d�����������X4��`	�[:X�Xb,�-,	�!�4K&!�q��Q�Q�P�QgZ�<fY�e�z�-��Q�G݃�����b9�
o�|��1*|����X*|��hmmuZ#��p��p��p��p��5+2\�H�h��A�
����V�"[�.A]���F�gQw��B݋z �����4�o�^D���	���7���bSP�6`AφfE�����555Ֆn˲M��=���~b[������I\XA�m�;Qw��C�FE�����cIl�~d������&ڷ	��G';� � {�o�`�b��Q�>�� 85�;�aG�d;�h���;�g��?f_n_c_o�b�n��찝}�� �19���~�w��?�_���T�����v>����O�Ok�N'8��XX�G�M�O��P�L|�|&��z>>��O�|������|V�g��g�ϳ>;|v��f>�OsW\Eu����Bb����Mi��"�EL!�0C@��F��4M��G04��R��Z�F��҈cDD��`jiơu�T(:e�ҔҔR��H��}���{��t2��/g�{w�9���{N�:u#�FB��Po!�[�B��z�zC���y�u����Ԟ��SPw
�NA�)�;u�LV�)YJ����+EJ��HY��(�*��'�e�ҬlR6+۔��[����]�}�C��rB9��U.�L��j��j����Uǫ��u�:K���U�bu�Z�V���
�qu��NmR7����]ݡ�Tw���ԃ�G�Q��zR=��S/j��)��%i#�Q�mZ�6I��2��Z���j��B�J[��i+�5Z�֨m�Z�6m�֡ui��nm��_;�֎i=Z�vF;�]҃z��鎞���G���	�d}���g�z�^�����z����ZBo�����&}��M߮����������?ԏ��'�S�Y����!��h���Xc��nL1���9�\��(6��F�Qk�07��&c��jl1ڍ�Nc���8h|d5�'���9�)�q�bZf�9�e�f����3Ӝm�yf�Yj.4���f���\c֛����l3��f��m�6����C�a��c��g���%+h�[��X��Hk�5Κ`M��YYV6cV.R>Rz���k��Z�z���k�j��Z�z���k��Z�z���k��Z{��-�^��:���<��)$�b��FK�ыm�b۰�;�k����)�t{�=Ǟk���|�Ү�k����Z{��do�[�-v����i�߱�����q��}�>g_t$'�Q�I���@���9��'ә��8yN�S�,t���N���Y��;����is�:N����v�:��C�a����:g��Υ�`B|���$$'�L���1\[xp'awU�N�]�vW�-�[�U��2#�ȵ��~ވ�����������s#~��_C�?,�]oy��5��v�������8�B~���@W�^����A�Q{�?�ҫ�Kt+���鱁A�{�����Ң�%���c�)�#i�cWz?�k]�컺��ܗW�~_��x�s�o���z+�i��q}��[�ף=|��G�GҔ���Y�pw�ײ{6}�v��a�_;7������S����>���H3K�:~<��_(<3�w��8:Ej�cyT'�W��V@8 �ƍ~fm�,6�Y5��]�ߞ���	|��	�!]�d�tm/�{}���^~_��t���-�e��m==�z�c�?�gR�}�ӻ�`N�o��) L�：�T��A���j+ç�g?C��WEZ�	�YB�0&~&���=�ITg�wW�p?���ȃ�wѷ��A�{=*��)�j��G���i�F��p�O>#�|�{�2jk��R�Z���m�u�[F'N�ʿ��9���T�v+a���}�^�#�pm�p�$���ϑ�����W��S��8�-;��mE/'F��%�(��~�c�L�a,�DL@.�\�3� \D��p5�j����6^'ǋ�	w�Jx*��%�+WD���3	�$<��_����=1(%�)��7�'"���7���#\L��;�_r�1v���pET��΃a���5>�� \A��s�N2��\�h�g>-?��2�d>`u�N�6�5��ؽ������e�]v��ҷ���9�{���ރ?��;>��J!>LR%�O�li
�,eH�y��)����~e`I��8��@�	<X��/ZyCLBL_34�V�T̪�U�M��?�R��ؙ|sl}l=9���'��������ئ�&��v^�_���v�u��w�n�v�-�!�Y>ƻB�C�y7�g,em1��2(Sk�����R(;k$�e�JYwPT���+v�>D:�$v	O �B:�t��iB"|��D�$S�N:��k>i:�@"vh���)qMH8'�J���.>�+D��Z$�Ԅ$"�[E,R��]Bډ����8�G;I��x����q��H�ٍ�N_B�Z��gy}oY~~�����V~��"���d%�1R�m&�S6���J��ճF���ƶ��źя����;̎�֋~t�]�A�5��d>�����>�O�Y<���|^���"����G�j�o��y3��7�m��;q������r��"~�K��ĿA,�3�&2	%ʸd�k���L��i�7)I�Y"�"�S�G�W��I���h�F�/*����G�/����܃��\�)����ٷ�,��y�o�g�}fQ�g)�}VQ�g�'��Z�gL8�2��)��O�j�����ِ~3A�b��w��rg<���̻������-�����Oy��:��B(/��d�~���c�L\I�~�{!����e�XFY��,���b�=�����TTU,gy�(a��K�*��E�p��
VU-j.��]<��h�>�r��Wz���uq����Y">l<�Ħ�Y�\ӅaI�XCÿ��N�c}�=�����(�Re��֕��
]'��*���!`��r�Ej�d��S�v~�g�f�]���L������Ov3�_�~���=X�ے����(�6�9��I��sSXv���������=,�	�l��l"�	S�.�f�=p/�߄o���](�y� *�!X�����������<����x	^�W�5�3���_�����	7A�@�����P�
�c�"�8�\�\�+ڡ��rshlh,�_$6��3�>x �߁�A,�e��~?�����Ix~	����"�������'���ȟ��bAS��`8|n�5X�1 X,B�,��V`bE�S�u����%_�4�~dA6�B@�BTC��
Xk`-4@#4A3�@+l�Q�._���=�I��|
�a(`ȗ 	R����g)�g�zЎ��Ip�_����?K����J��0v���a;�S��;��y��tҙ7��5)I�Q�E#������d�¶�$�	�j�Ο�и���`el�����wg���O��h�q��?N*3
endstream
endobj
20 0 obj
<<
/Filter /FlateDecode
/Length 430
>>
stream
H�\S�j�0��=����z5m�@}д�؛���Fq�����l1֎ff���z뺑�w�7;�й����i��Α(��1��mN�@E ��O[w�i���#l�G��c�����7߲�ܑf_�]���0����Hs�*j�z�����TD�����x�������TF,�����P7�kwdZ��S�r��ص��������},�մ��̟��V@����k ��S$J�B��@%�AX d%����O	��O�| A��Al�Vyh	B	!�!��(�7D�<�Z�v��eu
uu���M.dD.d�\��Lg��
�L���^L�&E�	��&Z�a�l�`�5dm�Y�Y��X4dmj|Z4|ڇ�Yv�s���Ş��65���00qH�L3�9����+�� s���
endstream
endobj
25 0 obj
<<
/Filter /FlateDecode
/Length 14451
/Length1 34804
/Type /Stream
>>
stream
x��}xTE�խ{o'�KH ��	y���!&!!�I���t�Ґ�cw�����0�ddEYt_�.��Yߢ�8�(�� 㸌�0����Խ��Dgv����?]ԹuOU�:�ԩS���ی3�z ��3cF���'�d��w��?��x�JMc����̊�?���[�C��U�
?���c׿zy��;�n��߃��뚼-�wL��X?�WNԭ�x/ydcC6���-˚�;i9c?F��y�-̅����Xָ�~��C�e��W7�����
}�Q?�����?lHCSd�O�����}�l�y�>tWc����M��-)��h�{�i�6��z�8���myK0�6��0�a�o	�[J/���.��NJ])��x�/]�}��	�>o>7�D�z���o��$T��]I�s5�@���M�I�7�R�G%�q���� ),�(��1�����<�4ƴ1�q;о�_�z�:�]�BWE��eYo�����QǊ�b�0�e�if��j�-e�}�}9������?b�b�]l�?���ql+���(�,��]Şfa��ճM�zv3����Yf52���o��na{�֊�C�	ףl>[����7��"��M°� c������v9kC�Eh��բ�&�}��D�u��`���^V�����Ͽf�c|��.��$K f/%U�����(����(� �A>��`ϲ�2���A�=Nz�IL�M��S��N	��Z�ޑ��/�r��j��T��@
;M�dS0��L���[��LT��VP�ϷX�3���.�:�1#��n�QP���o�P��P4[[ �C�6�� ٍ���iy݀���s��!��2} /�z��}�����F�Q���f�ǰ�6�r�c�X�Y�fC�GOi����K�`=Xz�(���(A�K���,��m��G,	�V��-�RX��J I��/��l�/���6l��i��m��>R�hK��tf-�B�b����r�i��6ǃ��厾��m[��2i�"�_4{���)9j�����A�����Hm?����Y�|�:��R��l���dZ�6#נ.��Bߔ�a	��b����$(܈��
�?a�(M��6�U�;�r�J��g��4zj���!Y�8ڂ4R��*��]�f���5�d1O%H7�yH�y��ߏ�>i�žd_*�|e>���=HT��7�>hW�q�7_���|6���#�X��� /�%ڐ��0b)�I�v'p}�/����ː��^��������W)����<��-Jh�F�ɾ�2>5�lN�)��g�׸���1�?��C�_@7[s?Oۄ�FY�g���5��<3ź�'K�{ pl���C��A����-��ZXS��0�P� ��>h&�R���fkqO^��>���H^+Y��Z�c)fv+f��W-r>ka�ia��ہ�'�ť� ,�ð��J
d���Jk|+x��9���=���c��z��W,�V���B�oZvCiR+v��1�b��l����ʐ���j���]����%h��~(��9�K��nl���e���d��@�c!��4����H��M�t���X$���]�a�u�|�P�F<m�{�.�~���0�_J�Mz�}r��٭��N>fOܾ�K~�!s��1���h5�ɳ3�X�$��D[��j�r[ G��t���|��9y0s1��d�A�������л +kOe��#B��(l�T�}������Y�n-V���<��.\w��C�����/��i�Kѧ��`9�9��)H��f����>���Rd�߆�#�s����g�KHS���G�G���b���6��06;�~�.Q�e�\�(�|
�E���Fhkf�>h�Zȗ��-�_\�G��c��h�}��?���ߌ�F�S��ϙ�{Z��uH�H��_=�e9��<lV"�8��۰�%� O��Y�_Y�lOE���A���C����(�甽��|j?��a����¨�z�9�&���]��pP�O���aG#�Iv�g�l^�4�O����}�.�<h�?�G�e���HC�r�s�xo>4ʑ3Q7��ep�Q35�Y-�+[��rx��7�4u�K�/D$���Z�2�i.�dB�����~&|{xȔk�b�h�FU]s|du +RFT��h���o�k֎���K,�R�q1�̴N�R��T\��h�l�$��$����!�B���8��g�>��/��e��M(���46�S�َ��<�K�n��}[�f�Js�Ume�'|�}�\�T+��˧�ooh/�Jx'�6�7�?�v����v�f�U%��?��1������C���<s^\t]k-F��ӿ6��O`vJ�U��O����\�d�X#d�K����:�;�Jܼ��%�R������"�w�#�S��f����_ �c璇L�y_�����؟QGz��V�p�	p��tІD����3�lG�Q8��1'"�(���
|��pV�3ըXG-�-�����d�ζs:�Mr������ �+�"��=�3#������/�v��y�+����$J��JP7��p�P?�L���h���\�!�{�=�By�N�p*b�<i�}P�f��`�-��g��6]�=y������M�#pF��pΎ)2�N�:y `_\Ӱw���;����HSXI\]a����$�3얔�D�'S!����'���Ր=�X��]���=H��j�N<h8 ǧB�+[^;S�֔aGY��g����΁�d�u-�հ+���p�L���L��8i��6N�w�g ���ѝ�҂Nw�"umAfٷ����l��D{y�L�{�3R^l��m�_�����j,�2;���4	3�'T�h�PV�Y7�h1v���Xm���n�~ʿ�>���DG�V���vf�sځ�|��,<�t��3v^@ǩ��z��nK�L���z���2�k�z�t�ڐ�C�%<�]�L������ S�o���Y3b�cJkvj�U� �_�z����)���JQ>�c|5�����g/���> q�@8�� �:��I	���:�Π��ɧ~��[$\)�늋]�	G���Tu>�O��NeJ��Z����26}I�Ys�B���H/�d�ݎ��N����܈]�N]�-�s�ގv���$�U&j�"����Q���Ъ_�{��������X/��}XS����'ơ�Xv1������څ����g�ଵ�����q�Y�V����<�B7��TB$��]���p�JSq(bC�S���<
+?|� ���r�Dg�6Dt┰'��ثfC����l��j9|���bv	�v�_�`������q���{�5�?�^ ������ �0��a�24ǃB.x%ow��]n�BgC�I:��!V��Κ�S���)F����T������������%��v���$���O�o ��^���ԇ�祈̣��V����BB����H�0�t��ѿ?D�Z1�# ��r�$�U����g�|8kG�B��vJ���W��Ѓ�_}��T�/��ۈK@ܝ�VoG�!�RyV(��]�o�	�vVT��8��8g*F�Z&�g��#��o��O!e#��b���®�e�����w�ZmV�\����s]q�]JgQ��Ʈ=�����Y�J��z��<叕��	w#���d��q�~��C�q�Wq���������?��m�:_��#ʧ5�<)�v��G�O!��+"=f�f���bՒ�s��ў�&�2H^f=��|f}����*���둨<�J����u3f��O�D��!������;��a/A�ɣ�>������%g_X���F�u|'!��`���~�8ۇ��,��d�7�O�0���l\m�
�e�)��X�sK�Y �5�մҲPkck��G]�ϻ�!�Փ�!�%5;�s���|��)ڨE���N&	�N�D9yr���W:y!��cr�?��w������>=5�?���m
%,F5kJ��+%$=��������tM
gٞ�������Kk</.4*�˭'����*�w[�9hY5j?m�~��~14a�:t��o�<:*{NE�g�3�E��E�UՠHw@_\$�h���P�+Y��S��5����oM�O�*��#�L��S�ɧ��O������xJ<1S<�'k��G|b�xx_O��b_O�PO�)��S7m�)�O�Ğn���b�3��j�.X���I��{�؝��$K�2��ybg/q߽3��Lq�A��|K���ڽ3ŏĎ�i;V�����vJ��[{�m�.Sl1��L����)ڦu��;Ҵ;����hw���S�m����ĭ��e�S�-��x�m�Sb�z�曆j7/7�77��]��������M\g���!O������'��)�i�|��*q(^�'֢��<�&C�b�O�2�JSD�ݴp7�2G���тږu"�!���ҚM�ԸDkzJ4�WC��%�1_]�B,���D �*Ч�'���'�1R�@�O>Sԙ���ub�).��ŗ�i�MqY�X�'��-L5�b�-0��<1��Un�:ET�E��Ze���"E�4]T��rS���iemb�O��b�)f���f����b�)1󔘱N�Ԋ׉��bz�(H��i�����Ŧ�:ŭMMS�b����61i�[��[LZ�Nt�����ڄ	b<��!ƍ����cǤic3Ę4�wQ�������;:#?]�-�3DP9Ũ�TmT1ꠒ���f��e���
�������b�A��F�Iڈd1� _��@>G�..�#��dhYC�P\��C��!bp��쟦e�A��ڠi��g���_�vA_1����&�D�4ѯoO�.�6վ}R��=E_��>	ݵ>���@�H��t�Ko�&��	�'��<%z�Ԕ<-��HAmJ��\�u_'�q�\#��L���pw׌���]$��2���"���	]�p�����%jz�����U-Qh9�mB(�41Pp���!�A��>�������c�`����`׵�q^����oQs!r��X5�`�;��Uj�4�� 2�E��L��QJ�A�sD5�Q\od����zY�IyY�İ5�4� �ڇ8}7NEO#V:���<��~�����\��I|�/co=��ؿp�wq��U��ŞgGٛ������|K��]�UlD�z�k0$�Sl>��,��Dl��!�^٦<�.��*�8�,V�R����R�����a���6�9�ڃ�,&���${]nsB��b�v���w{S{K��"p	.6�"��N%��v��|��Z�8z�)��	Baf�ڠ�B��b}�����VQ���G�]�R�;r,�g�ԡ�R5��tX�;�{�͕|�>4>{ŧЃMíAt_St5!��KG^�S_���AI|j�1�kKIq�|�ԫ@�`/�$&`�֒�����������NK�=�"��Nr)�%�sk��~�w����E(.��$��DE�C��R�u��N��ua棛9_�_�=�{b?�e�r�rI�%�7+땇]'������,����h1痉�q#_�o��͉�7����I��;J|��BHx2���d���ꚧH���O����~|P��T1X��ϗ>��5w��^�_�l:5R}�=���jW�����B�ݟ`�A��藤�sy�A����6���C4�
k�>RW�2�8Î�`t}EC�Ć^����a�=�2=�o� �./�4�q���OK9��c���Y�3�^i�c���i|L^��epfօ�0C���+������l�i��>�-�|�QF�<xp'�2~��5�c�3�Z�n0�����:��s������Io�n3֤4$�"B}{�l�>�/�D�~�����M�=,5��K�c�MP���[k�c�,.=P����M۶m�wwᤑ#�D��{�I#���س��I�I?����N1R?�o��&�6$�5$��o��[e�J^j�{� iZyyg�,u��TRSz��K璟qRm�7b�7���g����E��Qu�g������cy��s����_���:��4��J������zm���ֈnwfH5��Ό���~��������Î���|r<�d17����j�W�_��j?mILc�Xj�A9�NH=�Բ�#+�O�_��+�ٞȷ��x�I%��_�0b�79ރO3c�Xu�u�/�Ȫ�����&��7��֍���e$%lb�ueSRXn���$Wrʑ����z�x,|%�'T����w��7�Vx�y�_����U���p���C(�^۞k�� ��f�����zC/����^����9"��!g��B��\5L��Na�3��X�:�|���ͼ��y���_���;~��������w��ϛBz�_�8|<S��s2<?-9M$&�4ѐz��9�[b:s�J9r���>r8�6[�ɼYI/Z>��ks7�]r[VFO�|��GWM�#���e56��V��[П�:��U�Hہs�E�Z2"�M,�oNؔ��N��MO鑜F��^�&M"՞�
.R'I��MK��{a��K%=+��k�%�~}�Q�C�?;�玶�Sp��w�(��1+0�u)�Y ���jP��9UxΡ�`�9�M��"1�����qޤܘ7Mp���5:y�t��Ӕ$�	��"6O�S�	���Џ������|��T���^@�X���ME�#��wH�R�sY�(�N*�K�ez�rBL;�Χ��|:�Χ��|:�Χ��|:�Χ��|:�Χ��|:�Χ��|:��4��yr�O^��������e����)�+�W��3X�)�'[�X*��)�� ��)wK���㔓�XF�ρ���N%�pʜy�Ý���s��`#bx5���w�S�Y�;J'�e����l��1�ܭg���)'��cӃ-kB�eϰ�ូ��1��5��@$	��Mٞ��OAc���Z�=���?����I*�/��o��5x����o��	4{ZZku_��h����6�=s��AOa��7�
�͞��1�TOգ���Sl�p0���L=���֜p�5T����s���ѫ+��>�꜖��ѥ�:s�?C�&�H��<�aa��S�o�����$%ut�^�M9���Q��$%���t9 =����o�Vx��]�$%U�CM���.Z7�C~��,�m��}ٞ��G7�e{"A��y�����4/�(u`�ZF��Dx��M-hN"��hk�3,S�$s8��<�p8X�b<h������F���@#t<�(���`}dt�9\r򷄂��:�$�@�@mk�/y��!�T���#NV"���i
8Q���J�m�=���i�K�������Ȧ1GC�������ehbd[H�Gur�U��3;�4Է��1�_v�=�`�'�Z��_!���F�$	Tl�H��䤤jTyk�+�Rۊ$1#hF0aK���av�'���P�~Gk`F��$g�v�4C���퉬i��{1P��T��&�����dh��L��|Rr[u���!����Ɂ|�p`Y�dcY㚖�0u"�ցH�zD�	wɶ8��0oc�.D�~Q^:(����5�@'S�H!?��K��B��Is]"~؝�`U0�{2ck1�ƎVx2i�fJ�av�^���j+恄X��`�x�--Xb��F?U��r��i�F<�0(��;��uX���
i��ٯd��kf�p�X�r�h���F� X/ц-޺�ekn>�?��au
N,�뉩YŞ�e՞���
*�=%U�����%E�E�̂*�gf{�T�*�W�A�ʂ�ꅞ������9%eEٞ⚊��*Oy��dnEiI1p%e�K������_Yy���dnI5�V�ˮ���*"6��r�,����T/���(�.#�3@��SQPY]2}^iA��b^eEyU1h�lYIٌJ�R<�B���򊅕%3gUg�S5�ٞ�ʂ���s���r�\�Mr�%hx��S�Y������₹Ԗ�3��|.�h^YQAuIy�����ۼA��%s�=EsfWuB�q:�Af�W�f{�*���Pz,�,�^-[B��D�dwzyYU��@����Y�rP��%gR�2�Kt��+�c�,(�*��T�T3*��.�'z���O��2�_�#ihE���JA���8�-��xu��%B��,n�=JWj��li���	�l�µq�{�ʒ;���:m�َ�%���nd�_�J?�`�\	�G��ɪ@X�tl�MAg�{1z�Z�_z�-c��n�-� ��
"p&o+���Zg+9[UW	h�������T����59h��LrhF��.�W����2I����x��tDP���X�-c�=l�c�q�c�HcP�E+D�#��_�&�֌�9(�?b��������G���>�LbE(-���-���*�dK�D�*̀-�u+���Ý�6��u�S%���hՌL<�ׇ�AX�QZ��-�M�D!�?�{T�w�q�e�-]��I������+�>킸���_�IIs��"h�
\�@-����Q��-��J���3?�7vTO��:s~�.,�����44�ц����2���lk܋R<�g�[����4���6����=��+g�IjupA����B�UHzM�Z��ڴd�ߑk��YڣOҩ����h�۶�-�
J�e�g}�#A5��p@Z�-K���(͈���U����z���yo�d�4[�qV�)g�+�]Ò�:��:��6X�l�T"�&�z5U�c��b<v�@����`-�vN#v�0-�A��*����'%�H[��<Fdmt�o!�YKu�UR�u�J�@��G3M/Q�~��U�ܶJf�����|F�c���;��Ȏ�9Zz)��l��v��j��?��Q��ܶ�,:���:$Z%����F���z�a�	�q#�$�1��U����"�6�v��x���ɱ}����d�:��^�����s�:4p�'�}&⬆p��ѵ�rV��#e�:3U��Q[��a{r�9�3(w$�3�M���;f�ڬ���K/@�s:i�\}I'kb�7���k9�ш����l�ͩW�\�c��.�y埢��h�w�$�4_�q�X&_�G�p86Rԇz��ض��~��*S���u�0����qpnN:��U/g�1ۙ�F�/p�r<�_��ԉn�Yft�t�E����w��UR*��y�}13&w��>��f�Y��vJ��3�r��xmu�Ct&V�6p�QLq�j݂d�b^�Y����o�|�� =�G^��~iQ�l/�tg��T��D����<g���i��5v�e�#It�EWE��$���L�EZ�
�eΌ����w�?�'<�7KU묑��/��4E/��q�Y�h�r�U��'+e���#_L]�� �.F�y)�5T�)W���b�|A�ǡQ	H�C�=���}hQ�bV#�(�/������\`Kq-v�Qzm�<�Sy&�h�����ڡ~ċ�i5��v�D��l.�*A�S[ �%��-5E��3N���2ќ�J�a��Z�vUR�Rf��2)��۲K왰9��kƦ�R�j��T�̖�<E�?�:Gbm�ʝY�r�G�6�������BE����j97�������ܘ͓�H=��
ei��YkY7+ӥ�hވ�"9R��H�Y%�R�<;g���3�|�RS��u�X��%1�m�%R��nm����6Q���RF��K1j�cSRw���W��!�=�����/sfwzl�˥����r-�Vr��bZ�!��\��yq��y�}��8���:���.�æ��I{*u8��i���ھ��Z�<������;w|����ǟ٬���G��)�6uiׁ����gu�y�c���\�S��wD��������(>���8ݎñ���?���d�������`�l��qm�Z�]i��WF4Z�,�<�����"�{{�U�q"���iK��]Nš.��o���,ߦ����f��R�O�8tC,z>��	i��.��ˬwXQ�̺ơ��eq�����W�1��Y�c]#�l~�wM),�)���*�1��[
�΄r3��F�(mS��|��#�w�W1�^��̄�Q}����P~]}�7�P>���q�G�����q�� S�����Tf�C��Lb���L/�QZͲ�!o-˭[jdӖ��+XE�7�a���f(M��X�;�%E�/�$ƫ*���qg�3�
�J��z��9�J8���L���y6�jNA��C�5Y_	�$�iZѴ�Z`E�L����[=�/��r&�4֟�ԎeS�J�tIu�smF_���y��f�>q�}��S��{�Z���O�?K�d���+���>�Mn�=t�[�P�bsњ85�LP�t�^�ވ�P�U׫�K"�HC�K��K���e�-b9{�X�82-��������j�aV[��ֹ�P�+ۭ]1����M~��&������s�i�(\yɢ^�%2)�5���	���+�����^q�	�h}�?����?�0EW����T�(#�\e�2U)Tf)eJ��HY��+�JHY�\�ܠܪlVڔ��Ne��Oy\yRyF������;�c�s�K�k�PD�Hi����,�-��D1M�٢B��E�h�""֊��&q��"��b��+���i�xQ�"��w��qL|%N
SU�$5EMW����05G�NV��j�Z�֨��>u�ڢ�Ī�k�N�nu�z��[}H}T=�R���*[}O�P�L=��POi�W��C��jC�Z�6^��j��2�Z[�-��F-��֮�n�n�6km�vm��Gۧ=�=�=��R{I{C{G����������vZW�=YO���=K�����4�H��W����z�ޠ7�}��^�I�]ߢo�w����~����������~DW�@�D?����M��Jr���]�]��a��X�dW�k���U�q]�򹖻Z\+]WcΟ�N 6�R��R�i��MX�2ժ��V���vX��k\��ߥ6��=���?��i�f՚�%}��zkk*����`�O�OZ�\dv4�K�y�\ �6���*m	N>f^�����mX}�SX�����X'�̏�Ç�����c��i\e�5��X��]r�2�����/ay;��K����3Ⱍ|LE;��2�=�0���ܞ"G(k�?�Iʥ^f����.˄)�p��TKh�+��YB��0k�n+����O�`M�(����0B3�w��ն����}���k1�fs����4z\����r�������k�%1ci,�8T�K>��
�%�*߷�P~��_m����(î0�q9��N�+$<�܀�� _op�9-���(����q�g� ���h�%,1�4a��'T˿��YW5��.��?K�P�f^�Jv���� /��u�ϳV���[������s���u�5��	(1���%�/����"�~c]Km�M�^������.�@rn�/��_�*�_�ߌA�� hz���O3��-e�#�0庘���#��{�c��P��liC�\G�(��3�9��/���U��X�d�K�LҘ\�~�t��_ �H�Y"�qT��'�����:C����x0��Zhu�����,4����L��$�¤,��)n�Ive�9M���$���I�uB��d���������,4��,lL5��U�tĞ�����'�q���߳�;��+�l��]����U�S�:�33a@��ڿ�Ø��&��:�]�^�ޠވX��7o��nK��0���q���~+e>I�z�o	�u��3'�s�,Wi7hP��N����$�t�ο�_�ӊ�$(�J��W�(YJ���LT�)E�l�B��,Vj��Y�(k���M���e��C٥�U�+�����W�#ʻ��'�1�+�b
U$��.��L1L䈱b��3D��5�r��E�X)�׉��Nq��&���C�QqP�ů�k�m��P|&����T]5�j�:P��Ps���T�P������"u�Z�6�!u5,��Vu�ڦnWw�{�}����3�/՗�7�w�ߩ���_�_��5EKВ�4���Ѳ�l-O��Mӊ��Z�6_[��jZ���j뵛�۵-�Vm��K۫��hOk�i/j�hG�w��O�c�W�I��U=IO����z�>L�����|}�^�W�5��O_���+����������6�^}�����~P?������������O�\̥�WW�k�k�k�+�5�5�U��*sU�����]���k����[]�]m.�a]��&Ў�V���:��Ӯ�����
�W4ډ����|�Mܭ���7��]V�jح���<�'*|��'p
��t�Mc�*y��yKG��h=C:�R+����]C�u�B}�i:ED#���A���-(�Z)h�,�Z�R~.��b�P
�tI�<d�Vج<߅�8���� N���!��*)*y�b(���3�.��7J�/au�L��J�T��U��JU�H'kt���7�(N�L��T�F-3���i5�i�)گh�k8���I���K��]�$���`����?��7K�)u���v�^�H����mjJ����?�6���
«��R�����%�"�r�? k�e
տI��~A�d��8vJO�B>OCΞ�~.1'�Hju}b܎���Q������M��=��\�@��"�Á�L�f��(�zҒF�^�S��c�ƈB_iW#H.%GP��F�����d����P���Ү��F�̇4��C�g~\�:V�J�;Y}�P����\�t�#�W����}����u��K���tyd�X4��N��޴�$�f��Ȋ ��8Hq�\�O�C���tv!�x	st�HP��#��k�]ħ���*�$��u���W(���f�w�wO�t�����n�8�������f�J<��'4��Jq˟�f���[1G�H���Q4�4�i˙�1����dK:��
�`J5�@k��]�'�l9F���k���:�n�J-� ʂ,�q+0}��|���?i��9��7�>w��gHz���,�^����)u$�\ySR��w
9S�~�Q��R%]��f�<N'�x@�3`P�)m���<g�3�|��"�A-�EPCd5NFPW��UFPk�K�B��(Fu���>�q�W�Q��y�D�0��<���t��V�x�'�|>���J^�/�>�����j~����w�m�^��?���!~����������N�[ci�o��c��p��;$�צ�̙�g��ߡ�Y�K	�zT�+/�+Ƿ�&a^<�����~m<Wߥ,)���.�M�f$~������|.��~|쿠�x��\�Ņڗ(��X��,�K T`����'�XM�.;٠�@�ȑӜ� Wh���wr.��dNlel��5���4�k�c�e��4��O/�ey!/d���O����T�	��]��ĿbӰ�����)~�*8#��8saEV,���f�5�NV.�w3��O�d�\��ng�&�&�ܵ�u7[����5������{��A������,���~��ݏ��`���o�U�wek�M���
��Uz�^�72��ٿ�A�?�����X���&F�?��W��/��@ޅL��ݏ| �i��_D~�hc�e�����ѝd���t�1��#��k��|7A�-�kd�y@�� �+�{�}�>aǰ����~��Vp@��s�_�oj���K�����X��sV�7��.�o*Ǐu��
���/˧[�|���s?�1z�n�l�>]g�ܱi�诓˿L��T�[;[$���?;�9p��ߵ|}��/���1O>k�!�5��g���Ycc�SÎ�����%��u~樝��$c3�{zA��UWU �,(�O k����F>���O k��Z��F>���=��1�lgz��db�7�g}��elZ}��ˊ́���U4��|	7�}V��,���;�,�q�E�.iw���P;��L��,�Z*�z����w�+_$U'|�z�Ko�S�h\���(=�Lb��Cz���lA��� N�f��F�1Øm�F�1�Xd\n��F���h4�����Xk\c\g�d�j�il1ڌm�c����k<d�s�r������k�q#�Ѝd���a��M��1�b�02����D�La�#������\����2�ڨ1K��bD�����z�c�q��ٸ��jl7�5v{�a�~�i�	�g�c��/�H0R�4������[a	�bD�L�\�ֻgdE�}ź�k�G:���e��ӷ�3��F����̸¨3�F�Xe\e\k\o�l�fl2�2~`�c�ظ�x���x��7��?u������2�=ݖ�ϸ�j�����l���4� �gL1f��A��`���CP�!����Ҍ'PSd<�o<8-Vs@�<.k�5T�J˕߄��3`�� K�Ŗ�d0a���J������Ǌ�y�❯���熧���)�X�	`
endstream
endobj
28 0 obj
<<
/Filter /FlateDecode
/Length 265
>>
stream
H�\��j�0�_E��Eq��B��B.v`����̰��q.��������,�B�Y�=wZy`�Έ=�JK��Y�@pR�H%�N�3������s�Gu�#�68\��؛�蔞���������Q{8AӀ�1z����,Ɏ�q�c��e|n!K|��0�:�'��������_�B�a����<k�+n��Er%=�%�#���-х�$(�JA)�^�"ʉHP������g\�}	bu.̟v��#+��o��FU:� ���h
endstream
endobj
29 0 obj
<<
/Filter /FlateDecode
/Length 2784
>>
stream
H��WM�ܸ������I��D�00�����܌�6p� >l��!,��a�U[*�)0ƭ��y��X���h5�/:����&�2y��{���ż���������S����G3*������ˏ�o����'���U�?�/?.��f58�������\���F�1��#<[���.~�������+�-|ߍ�;���:��;?���������m0ʺǝ?(�O���Z8�UaHǾ����|��|�:���VE�/_�_?y�#jH�������yI�L������@a���5�ݥ�U����� i0�\��kzV��>������~qRs�L�<\�Ň �x��;N�؈?:5ω@~ڨ����J�?6�iw����H	�M޼��`��,�a�ez�'�j����j�<��]�S^(y���ᇼ����"�Q��&߷F-�0)�օv��x��� �8�]Kl|;��@ ?�Ȁ���ѷ/�0�b*�k��b��l�W
��WJ�;ٴ*�$��U��XFǂ�b��D24�*_g���Vˢ����K�}�&���hL�ߘX�k��H+_`����������k-hg&�S��v>��>���g}@��s���4$gjgJ�G�8��� �8�ƌ��	� ���{F��|��h�#�?�� B�iZ<�f	�8���kc� KFC_Ol�S#F`*ݸT�,q��.�s�xt,��sP^<�SϘ1��g���
��O��
{%���iz?(�n� �c�������F`h<b��M�pI�b������w�͝�Y��t�ol�Z����Q
�ZQ�e϶�ܫdd�:w�����d�����ޙ� �10@���a>_���x���kՠ�\�*������V��>~,� D����\ư����[�#X�k�q��`�=X
���M�K�&F3���ތc��V��/��I�X�r��9�m	@��(>���i:e�>�p�zF*a�:�<�+V��k"a���t�s���^�dN����ޒ��К%�"�x`Ot@�u�n8D.�b�O���X1�{�N����5(�S6�
lM"������QI�o�Yq��2��dH�2X������{��t��k���21�6�w��ҭ;�2�9��ֶX��Zo�[C4�-n�z��dۘ`,R�����,�}�i���"�s1-�^�[<�Yb!~�X��=#�0I����i�
u�U��鸾3���4�����t���9X�
*�6tE\��#��|���ӣ�o4&�rV���_�՘���ql4��D'=�;�:�M=��z��O��D�Xl���i�HK���$��68`�H��x��l��x�k�8&��Y�8�#c��@: (��qu����'�֜��<r�1�ʮα��^��	|)��O{{!��jj�����5�;/������m���R�6s��KE����P�Y�9�&�YO�6!�5Q�-e�o8X"ޗ;�+��L����']�$����9 ѐ��+����C�N�кs\��lĥ9v�ȶ��8	Y�A2j���6`��K;@e����:����|b<�J��}uT���e6��fz�=�5��0�^�s�u1�����Q�b��W/�����lg�"�Q��L���) jMA�k���0�pM����{���jf����}�e����o�4}t��̻�V��l�JF;B+��Y�`���!�v&���U�&��L"7��y��B�OtbwN3�40�/a		^��\G^I�T�Q#?-�6p�}!~�TS
#~_�Y\�Z#t/	��TbJ��)������������2,X�'u��t:�3����NW��:����H����΋H�q��M|cj,����VS�;�|�)�}%fa�ʷ�۩��'UXE
�'NY����wX�-w����o*X��D/Q"�2����;�����^`;�;�[!�NI�;Kިo��*p�E*�s��r�x%eJ~㌿p�<ĉ��S�����`�AD���:�;i�7V�ddpK���ͪ��*�_"��w�@�P<�����JL�Ah��#�􎙵�1u�8D�)46!������Qb��x�m��z�كvwmq�$}hy�km5�B&�Q���JR�������!�v&���U�&��L"p�"%Ƥ��X�i��{N�%$�ic�mp8�Eb RU�[m/m�b�)��;C�N��l��w���ݠL}Q	��р�;�� l��ޓM�E��l;1i~_��0�䓶��U�5A�ﭷ�O�L��$�E�]!~�L0j�]`��nS���A���a���ΡHm�;���呏;��w�����y;���!Z��@W��ykY�[�n�z�5a
�ZS�^�8t/k53~��V)��ܲF�gǲ&�p��� ��h��w�	�]���2
">�5����B8��3�q��QI���=|M�C���a2*4�K��1Vg�eꬤE|��{o[��e!lg��Zu^��h�y[6���-��IwV���-�wV`��</�Bo}[�����^b���o�eN�%?�;���W��2����3�1�a��2t���§���@Њ���=Π��V��ʸ�u^r��N��W��2h}s� <Ԉ�B��;�z�q3zT"��O,4����A�B�4��2j_����R�P}�^L���d
�K�=�� $9�8�C0���:_�& G�x)jrqV]��7]�4��p)��`��� ����U&'<�Wr&:M�NΥnK�p!��/{2ݥaWs��"ƢbDĔ�3�1��`��,���_ ��o
endstream
endobj
3 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 4 0 R
/C2_0 13 0 R
/C2_1 21 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents 29 0 R
/Parent 2 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [3 0 R]
/Count 1
>>
endobj
33 0 obj
<<
/Count 1
/First 30 0 R
/Last 30 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/Outlines 33 0 R
>>
endobj
32 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227163233Z)
>>
endobj
8 0 obj
<<
/Type /ObjStm
/N 19
/First 141
/Filter /FlateDecode
/Length 2610
>>
stream
x��Zko���_1m�� R]�nc7�ܺ����:dQ�h���=��]r��Ҳ�h�9��ݙ�;w�kfT�5ͤf�	��d���DT)�:�j�֌˦D[���=�:8�)�;㽩����7>��5>����hд&������:?�����o�����ыw���j���l�����ns��<:}��y�'�on�����ٓ'����-��f�?�xz��g1��sq�|�z�����f�Kmz��͟]-�ߙb}�9;[��\��f�-�\#�����VW����z��6?ܮw/VW�`����ɫŇ�����ӳ���G������Vۜon���������ŕ>|��Br�����j��������o��i*�ןn0:�s2����c���e�����n�f�X��>�a���^��sx��#������?o�tf2���l��\Xs��Xzϕ���j%A��&�� �hRe�j�K5��|lO��e֡@MS0�9<�&g�s2)���;�w���	��K0)T���z���:�Ս%��
� �6�V�
�`9���NW��&04��c�ɳN�7̙|��G�1�g�V�Wⷡ�	�d�,cS.�+�����bZY@���"KȽ��c�^^���Lh�'�ȊH�O �h���=y÷��~���l�ج¦�)}���#6�IP����C_��%
9:]d��/p`%w��=��`�(�t����^��X/Jr٩� ��+�TQ�DY:��b�J2��a����@%��!
�)I�w������!p������1��ߎ2�A�Y�T�K���c`L�s�B�6%a8�J��9�V�ae*ԴP��-/�E8)P�Rn,�Z4C�RL����W,8�HdCh;*M�6�WL���^��:� ���-hy"D��X�lY��L��*RBċb�*���7Kj�|Y򘩨/9��ʨ����<B�����s.Y�B�e�X����4*5�#^��u�EBt ��3U�<���`��s�;1�;Z�m��p�0��A��c�o>�p�l����	�KM���Y�MAO�B���
7�U�+.U�/�`>rF�=ErP����uy,���eU4��s��װ8�1��ET�߀n�RO�����	� W�[/�`�Ȱbܯw���5*�0�$��F�=ư>�1�`c�T쬊`L�дtZ+����%���Uqb��>*_�Ah�Cy��#Cls�$O��[��1C�r�!�᪉���%y�Ԛ�ls�-f.4�6�u����ח?À'��m�>S�G�5�6��~�˨�(n�]�D;�ЃY�-�f`}v�ʆ��. �76����I�� ���uKg&@=̐�(�E���a��Z��]���=�������֜G�Wu��ms'�4c��G��փٯ�Rs�+5= �]�W�Z[�݉$[�;�W�e��M,�֛�]z�Ͷ�PZ2ܮxBZ#�[��#ɦ]�e�1�ށ}�Vۗ�D�	d�9�w�k�y�	���?�q������G��r����7��l�$;��z�]�x5�d�2vA9�=�
cUi��n�m)J^
��D�a�܇ZQ��q�또1
�՘�I2��a�]�����C.ݶ��diI�J��L$��'��&�E.�ߔ��J��jS��@v9��T5���3��G!�< �}�w�phW5�q
���|��g�o���C�zȸS2�B��N�E� �v_C
�R�Ζ��t��):��M�q��/��;���8�OT�& �G!0))�-�)�����%GPLT8Ǩ���c��"�AP�1��D��.sk��b-��^&�Ab�%H&2���ˉ Mn��1he�|�&1�;^�xW��b?�<�`����+�֒g���C,��
��l��
�Xy���M2b�˘���Ǿ�nx~FDqD���N�q8ā����N�����5�i%��c��G<!N�L��3���@SNJ��}�Y�8�l��|	�C8�=��2�>�<�%��`��=�}e����w<��:}�O����kj�!�v��c�:�om�>LBe�,�;Et��<W!��LRE�2���5��;T���Pw���*����_�7U��[��|���˳C�`z+�nq�a�;������o��x#9�o$O����{��?�Wh�4P�7�	3�����℁򄧶$���3�$��B�M���q�E��"Tc!�#-��cJ�P�E��"Tb���J�N��"Tc!Ńe�9�7��*�P�V���ڃy���\(���Q^��D�&H!����R�F
�Bw��cJ�P<�R�9�R��*ō�R<���`H))B1R*��Y���R�E��"kʛm����֙�X3���o����x1�t��v��EU����K�����9y����ӗ����߻�޲��w����Z*}�Z����8��E�G��Ù���vwd^�pN��Ŵ_L;��~������_k��>��;ު�@wJ�S�^�&U�?\��Q��~�R�(�C��q�R>M���P)����W��=���}��̿[�^C�B$�׫�s8�|����a��`b��?=C,5�g��_o��s.]�
endstream
endobj
34 0 obj
<<
/Size 35
/Root 1 0 R
/Info 32 0 R
/ID [<51888BEFF55B2B4F9AE414499E1C2ADE> <B6674D4A1CB375B00F582F65DDBCCAF3>]
/Type /XRef
/W [1 2 2]
/Filter /FlateDecode
/Index [0 35]
/Length 119
>>
stream
x�%�1�@ЙE]�>��SX;�@�9�&lE�	L,��Ͳ�߼df����p���
D&� ��u���o�E��(N�6���j�^���{��*j�C::mֵ����y��<�&�q
endstream
endobj
startxref
47457
%%EOF
