%PDF-1.7
%����
10 0 obj
<<
/Filter /FlateDecode
/Length 23
>>
stream
H�:��� �����pn@� 3
endstream
endobj
11 0 obj
<<
/Filter /FlateDecode
/Length 2818
/Subtype /CIDFontType0C
>>
stream
H�|TyPY���+fh������JTtaF]AG�@���G9�
����@ @ 9"�C� � �*�
�Q�x �%�:�ʪ�[N�v�-���g��j�������������ǁ�@gy�����u��D&��և�SU��rGq��+*\	z%��hM������
���ޯ��K�h�i?W�KĮ�U���z�q��ɒ��Db�R���ek��4%�����ˁ���ى[��͉�^�fooo'nv�ʩEEhJq���'M�ɳe�D�X����̤��
J.V�幎��ġ$
J,Q���T"[L���r��R�E�Dy%sT����+J"�X-*J*q�%����������,SI�r�X�a�ވHM���D��.;(-���\h-@�(��CP�p��!(��ul��e�2�dàph���wY��w3��E+�xB>���� V�3�Ղ��Km���9,z\���e�B��
�i�w��dj����G��P�p�N�8�`��,
M�1��w����O�;s�E�:/]ſ��m��5R^us��G�\�)e���/��'u��!u5�r�ᘾ���������X��\T��S ����'�ȓ02������,hmm8݃=�����L�p�'��s`���ʺ���� �oᯐyZ ~C�ךf��pja�Lh؅3u|dF�����x����@�@<s���
9�7p����c���&��Ҁ�����l"Lu֪Ny1>$p��ƅ�OGG��<�t�cu@�_9y �u���B;���~å{�5�Q��8�Ÿ�� x=��g �qt���1�.�/��Z?��ÐL
�	�0��ɩ�m5�dK_���4V���s�<��^r��c��ӆگ�b���Α%����U��}rzb�)pŞ�ݍ%&���g\<��������V=�ߚ�J/����7{`̖�ń��> ��+�e�}4�;G;�� ������y�|� G%���M;ѐGj,��o06��ư�B��H)?��L�	_��ޓ'��S]��FҢ�S�{�?2^)�݉-��~�P_k܄-|��y�	$WF���3m�M}lpCa?��?;�J����(S���c�08Q�U�%�L�g�|�v���"�Y?� �v��&�Ͳ����5;��8�bxL!�0+A��#k������l?6OVU�0�4��n�38�Ms���R�PZT���5M�Hp+���C����Yxx�~�L-�+*.)Ĕ6uKc}MsQ{�l�XuM�m��sI�I��d���y9�q��?���wt��Q�o*�	J�ۏ5�G�4i�9����1��u��l�mo�c����Q��Y.�.z�p��(�5ȷWo���zI���X��[���Fsq=i)H�$㢐��h2(:=h'F���'�	���{+ao��h�D��j�󿂢�N7^A3*y)U��1�~�F�
x��ڸCژU0b�UJ+�pf#d8�_L��m�2�$����Èl����Z%@���IT�H-H�L�%�������i�0�My�pf@�.��*I$��V��`I���T������{t�7:*�p�tD~h/��� �3wZf~ �`�z���r��`���"�#🛆�Fp�������?�z���֕@e�y�j����'[���G���_):�ޏ"o�TC�!� y��,M7K��?���Ky$��h�:#'����2�\h��T�K��Q�Z-(,<����O|�pq�,~���_[0��>��Z��Ѵ�56�4����-�S��/c ���ɳ�׍<����f37;��%������E��r2B|�����aҺ��~C=��N�G{J.������.���u��	�g�XM���I���;�o��>�z���t�c���UYe�
UVv���F��P|��7���K8A_�c��Fi�W���D,��*B��j�73 ~��ۖ��0SY�����]�����<_U�.��	�x��Jx��d<�1�𾲲@=��lp����"�@�z;/�:��%���z]��Ѯ��>��3P���t��,���1�G�-����4�7 �1�5�.���j�,�	�X]M9T������$�����?׎w����I����[v_Z�uă��I�cI��M�q�z�>������Ká������|�ȑ�����������s�i[`SYm ��!������������ƃ��vp�b/OPE>�j�o�t�s_aiofO^��yq�g�G�}|��x�����X�@�^�c��������cP��=������������}t�rrj�������������}�JIB]pn�����<�cʔ������v�;���0�\��q�I�FrĄ��|[uJk0h8n�c�q�{�������ar�����Q���������)���֦ǔ����������!��6��A�5�!��o�N��f�)�(������ԯ���Ȓ��Jr����ykyjwlwnP�y�������\r���Z��n^pcoh�cY��M�q�O�W�������������	�p��`�q|��v�1���3�V��r�I�Iră��evL`�
oG0��~�������_r�~�T�D�����z�~�|�~�vxht_wrlwz���{s�s������������4��9�ޤ��Ĕ��� 
�&�s|��I����%���������F�_	��
��w�n �U-
endstream
endobj
12 0 obj
<<
/Filter /FlateDecode
/Length 293
>>
stream
H�\�_k�0 ��|�{lJ�j]A��M�a����t�C�~��\�`��w�3~��k��;��JK��X���4��J���[��a�7��p�u?�� �郳�+�.r�p����h�`w�6{��b���DP� �����x(;��Ǖ[��/�k5IpL?#&��i�VȊȯ�ʯ�����qJe]/�[�c�EITnJ�AiBJI� �q�)&e��t"e�'RN��Τ���E��D�s�Q��:d9�D�=�s8��4�q���c�b�֏1\]��69��q�f2૶��
0 x��
endstream
endobj
17 0 obj
<<
/Filter /FlateDecode
/Length 23108
/Length1 50364
/Type /Stream
>>
stream
x��	\TG�(\۽�7��\��q'.���PqYe��Qc��D#j�H��8���F�[ԘDM2fO�L��$�q��Nս�e�{��}���c�[�nթ�թS�-�0B�C������߾���hm;8>!q��e-n����fDخ���+��38cDܸ� t�"�O�Vկ8���G�g�y1o�*B�ș^i�Q�X��B$2�lJ�X2�3�l6�gJ6̥ �žpo�R4+���;ý�_A^v�bG����^�`�%���}���ʙI�d���ԢҜ쮞=ap�[�=��c��5�_l%��y�_���Pn-��/+���/Dcz�.^V�W��	�o��6BWdB-�JZ2ѭ�O(���뽓]�:�?�h��1C_����S��v���?��{I�%��-.�P$�� +��)H�`^A�]��-ݥ�p�]�(�x� �l�F�;
�����3�#�����b��n��T/�E)�_MB�3�gb�˨@��BN�ُ�@ԗX�n<�DYx=��7P>Z��Mh9��B}%Z���x=�p�A!�%�8�x���<*�	�U�Z#W��qy@�����Ǡ! �P}�Bs N�r Fu���:��r<]�yO!n�d��M�	h����g+�[(Z����+��C_�w�ZN�����J�y~���:�����!�6��zB��Q�	:�Rp8��r!��@�t( �
���ƲZ��r�c�r�%�E��P�<hY�v{=��0��8������F�g��N�����ւ�b���o*`G�cT�+DȻ��(��c/��a�Z���� t���	�Y�B��-��(���i'���uO��\+����7�cD�P���T[Z�C�דh��/�A��?���A��n�;k�k��vX��:�}0�c��jGt�8�-�B��Yڜ��
�������i���V�k�M��A�Bw�V�U��a�y�5��9��V��� ��E�>h?����Os�\���,h���R 0�^����	h7�M �x*p_���9L�.L�AnP�A�/��B�j0]�y{��ZB�����^7�����k��t-�{�|�7<�#Ag��p0��D�����Y � ��x� ��;p �R��!P�=`L��{x5��� �"1f���n��� W��0�Gb���"�����d�5�w�!1n5��f/�2��9cexe�Հ#�F�=VB|B�{F�^ ��܇���U-D�b�o ��7��w� �_�2�۸��� >>������"W�x<S�`xQ���PO����ݡVkg9�o���P<�*�vhM���#�6虌F�=Ũ�b�F���� X�}au��V�g!�#4	=	�7Z9���l;�y�[	��G#�R���c�?��]l�A�T $�)���n���ŀ�C:���8�.��!z���Έ8�+f��1�����|�������}�B}P�{�/��$Ɵ��t@�I&�4N�^6���� �� ���f��! MF�U"`�4N�o���{�	n���,�h�}�(��uz+[D蕂�&�9?������_3���I�P�[�a<���,h"\GB��2	Z&�I�Y �q=�/�wz�ae��g�/�,��Q���$����@=�G�`1�Q��<ۆ
`@�}� #v����� z�����wG4�a��0V����������P2?b��)�=�}c���j���L<"����4=R|
���u���.�8X�AK�"��8�vt��ٟ�Y�@�5K�yH̆��c�>���h *B� ����Q����T4LD��< +<Ʌ��3^`����y�C�Y��ĺ�(�~����&�$�-��=;boq}N��M�9��coq�[�xF?��O�Am�^[	ϦA{	��������`�e�%�ԣ�po�d�0V� 14��� �!�c�c�uhK ���tH��p��cad�hh��";��!i��`4GC,��gY�a�(����� �ì1��0*D�
Zc�L<]�6��ܡ���h�ĳGqdU�2O�:gV7��#�r/��r�f�+V+4ϥ@�ō�e6�Ŭc�h�/�E��l�AU_�"���c/</h�g���@H�q:�
Gq�Mxf�\��<�r.ZF��� �Z��������"���>�>�ae�J��p�1��>�>�!`G�:5Ǵ���p�	;h���a��U�:e���t�ϩ+ J5��LP}[�	c�ŘW�?��z�b��d���b�K�MC��5w3����B�������������w��M ��8����q{ <�5�� �r��B1���W��N�-v��FC!�����n��{η"[��t�����T��Bt<�@�����Ga��U��MqR�-0.	j�@Tn+�C�Xh��p~� &"Q7���y\y�Qy�h�TWX�ҝ�-p����{�#�x&a�u�
|=e�����O��p�׎Y?96�龖8ܶ���0������1�=58q�Q�(h��<%���p��bD��Z�3]Q�ա��3��~�c3�{܏-��޼���ȉ������B�'t|O��
~��N�<��aO�=N�;tX���3�Q��,��(���0�Y}(@��	���è�Z� ������Q� �z���rd[1�߀� �~�~r�1:Y���O����k��\x����2��N4e����B0d�>|F�sWF�_�YunQGk���fw�w �^'�6�]y������x�ĚD�om�����Jף��}��;�O�����X�;� �3'�����_|r�~�W��1>ǟk}|� G��*p�a��3�:�t�����@|u�� �qo�
]��:�B-���X"�s~"�� p�B&ܲ���Km�HU�y�cv�34{>��_�O?φ|zԂ��� ������AD��"���!?3@�#��i��>�C�pp��΋2PH��,�zr:h�T�@�6b7�r���S ް����!�;_�Um�T�h� ^�����z-���:7�ـ����t�
��dh�k7��ao���A�/�>&��=����N	� S�
�]8�������
�T�NM���@���P� W�8�=����*���`ۮ�B�<-�`�B8�-�L x�{۳pVY��@�-�U�m��A	��J8�6
����QЯ5�"A��0O �[�������� O�!*�mE�.�~��O�{�%�!���[���%��ǣw�Bo�� ~p2�@��t�����8Mg�^�N��Q=���`��?q����w�<'Tp�yBo��
w����gF��ĻA�`�Q-�ͯ��y���k��#��TqRH���1�x+�<�1N�a�
�8�t� yL	� Ѓ�ca�
�?�|��㿆�s9X'���b��Ϋ��}��U�d�
g�I� �}�hw\{ٯjG��~��b���B�xTq�A��2
?�#�2�:�O�8��ɍ�~�~���_��|�۫
�W�z��
�W��l���ڨ� �w�j�?/��@r~}v���U\A.�C�F{ʰQi"zYd��W:�N�ŧ&��'%���#Ȥ?���,���w'	�Y����0��p��s�y�w���π]����u��c��0��u�O��?�
98BW�O��QhŢ�����C!�0�O�A���C�2V�pX�# �ND����,��gb�Cޯ#ĄX��I0{��/���r��v�W�'�_��	�/�,}�}a΃V��Az�r�O�:A1C�
���k����!�k<��P�9$I/a�z���sA ?��@:��2Z/��5Q���P�]��T(%Pʠ<
��,��3Q`�@?����/��I�ܧ,>n�/�~�����>/��C�wР'�3o�?|`�����D�v����W{q
� ��\��Md#͞�{�V����l\#�৉��!�ߡ��&�'\'��v�nG规Ѱ�Ǣq�����K�W�Aw��WYb��0�u?	I���h������a-nmVŶ��w�e���ӲXi�~��~b��B�����_t��e��>	�:لI�И�U~�О/��Y�K!�/i�~[N�m�uEp�
k^t�W��}`�x)�-��͚^��B*�=� ��]ԭ��-�]E���?K�!��-�f�!I��$�E/$s+�.�>��3�NE-8f�JU�6̣�*�Y���迏л������`w~-�YE�,`?��~M�a�C�?DH?ޣ?D����J���7��wi�X�ҺZ��;��`��\�ۍ�F.�F�����w�~݆�M�קѯT�����~����~����S�~�ҏ?�>V�G���F���������f�Co��<�~4�
7W������IzO���e�^R�;+ܥw�ҷ[ѷTzq#}se���J/���<zN�o���J�lq�N���JO��u�� z'��q=���J_;:^z�}m;z$D::��aGB�a����֮��^Q�!��G�����\z ���J�{�}*ݫ�4�?�t�J��Aw���]�ҋQt�+}a���BG�ӝ�ώ���̣;��?�t�J�Wi�6?�&�n{�*m��Y�Lt�J��I�U��yS��Y���i5�_��n|戴Q�πo=s�>��mX"mO7İ�*}Z�O��SG����6��i�x��f�
V�ҕ���!t�;]��e*]��%�ݥ%*]�N�T�"�>�'=�A�t�L:��y�|�>>���sU:Ǖ�V��NWiU�E�r�U��\c�Zy�UxЊV���TZ��Ғ�t#-)�(�d�⎴H�Ӣ�T�Fт{t����<��4g�������*M���*��҉*�0�,Mp��s�st,܌��c�<:ˋ�R�H��h�'����*�Pi�J�G�T��EST:w���4�֑M���I�<�$_:$�W���p78�&�]���K�!�7�.�jIL���źIq�4�� ���q�b�hl->w1-R�+����n��(�Ё�8&&�Pi`��=�O��t��*�
�K�tk-�F{��WW/��J{�="[K=���p��(���n�[kٚF@-�[I�Gh�0O���ZK��aVw)̓�qv7�.�C�.*�=;��N$Z�Ҏ*��P7�*N
I���h�J��ܤ �ںJ��+F�af��Si[�m[�����U�R_�� �D�ʻ��*�z{Y%���J=������*u���f��S��;7W���F�4ݹ��$Wu�t��s1Q��Af1R���̬RHbR��5X��RH�*��(��=��J$�b` w��Jq-�]�w��煺���j�P-d����O�5�d>�l��0x��_-~/Ǉ���^�~�&�����,�k�t�G��GU�(z�-A��/���=�?j˛f��3�S���c4N�h�����h>�+I�o�o���)�z��B�s������m��܀�� �{� ?*l�b|���d7�O��w���/��PC�����*�T�MF[���&��^�n���ɵ��Rp���Gq7�������L:�>F?Y0�Ao���Ip�G�*{��J0Z+��Yl��9\>2�M»��9�ޅ�@�].1BI��"�����I�հlEo�{�������D:��a�=��g���KiO��͑Vk�vt�VӍ@_hw'p�#�x%p{�YJ�Qo���t-��o��C��x._�nd���pT�Q�^��AZg���W�!땺+u����!���W�6�S7*�w(���,�NwSЭ��B8^��2bDf� $>�n������������JW�N� �w�?�*����7y+z��EA�CF�&W U�޷/P����2����	%={x��U�-Z\S�aC��q]}�뿩�_�ħ>�����n]��U�ـ|�����E5�����ۋ(��<z� x��Y�e�:��g_����g�����Y���h1Y2�B5�aĬWN�E�@�@�K��"�v@��������!���v�/�$�O��o���n�;�����q��Хo���e�#�O��W�i���c�7�KW�]=ۿb���f8UcSLk�?F�jK��F�����ȁ�M��`@{�Xo���z�fd����+A#X�!G(�c�)�<��@:�������Ɓ���T��SI�)�<M��D�D�6�o#��6�M�&oS��������}x�G��}�>y��ϰϸϴ�|���qz����Ǖ�������_bF��Nd���De�a��O�K�ڏ��q�^ݣZy{��A��A����=���J:,Z�W�{�IK��g���+W�^�r������o�&7{���L��������ĽpoY��T�O�3�2�8�/�q�a%"��3��/Z�H��LA�FC��O�2f0��za���|a���z�tw��⊣ս8��Un7�J�z��n$�n��`߶�јN�m�$K�~��O�Y���/�T{md�� ��`��O���og���N�p��Ox�b$�����O_~�s��z�={��J��{�)�W���UG�o����ƞ+��F�G�<:���ݻw���fW��[7�b���M:Q˿~���?�~;����g��i�q�K��Ҷ�mu�Fy����Zy"���j��A^ƀN�/0|�����z��f�H쏽�X�CO`�����*͘���[��4��)�g'�<p`Ӗ-+�>�d���Y�%]��r��g��Gh��={l\��杳�+�t�x�f��/sv�x��OV
v$5�b�uA���!jV�%L��ń�Lv��w���_�����:�y����΃�Ϗ2�@�ݽ�7|�=�gj'�A�o�q�a�Ԯ�����;ԭ8�8��Z�]W���Ĕv�����5^�.�-s٬���������5���������RO�`Ww��텚)���r��t�Qa�`��տf�Iw8���y��-࿻է�n��o��[6�[Q��o�9�p�_��V��M�Vӟl;kXu����!A�(�%H��bπn��i���������|�qy���RD�Q�p����Jc�~6p��g#w�|���O��p0��A�d��,[&<�A�L�{�4�_?����U�)<�h(:�c����w�X?+��<�ʨg��B(�!Lbqh�Jp��A(@^O�� �v�c��2:t	S��{�}�zJWG�[(u��v-�����"Р�_�� W�w�������H_K������݌��m���[`@$��N؍k�����/��I!�,���k�=�x::�1I����,^����§~�t���nܦ�ׯ��m�̚�`��Yș�+6W�Z�)3����/�00�ܶ׿:_sO����3g/X���|�)Q��=�)��V������V��m7m�)2�[B����ׁ��
��O��A*���ݕ�6��6n�P��p�z0��/���Dpk��)f?����H�@6:Lٰ̍�_�4l��OlTW���R�"�� b�eD�&ƅlG{�vY���V%����]�t��Y���Wl�@c���hHȈBb<�e�G�]�c���J;��E.h=
Լi�'���ԟْ�;y�;�B<���^澗�V�Yl�^`���F�+�Y�ud��Eq�߮��i$޸'f������?c��u��z��}'��풅'�Yt�.���Ȥ$��x:�1_�k
���ϟ��[�6���LhSL,
���
��E�$f�&b�&�/5A�S��~}�Ѡ��MC�a2[?���:�(��b�(�?�����b<>��	��o|3�̈́Q3*�a	^N��xLE�H�I�U�_�	��\��S�e)��ѽ�������v�<��<�l<*��j���c�6��n��4	������v3"��@�t}��N�4������JH�����c����ܮ������ԡ����.Z�����o5��o�d�꧗�|u@ټ�rw�����Z�S��;����g��g�o�ڸU���ͨ�(K7���|��<Wc
�5������iC�Z:aw|�/���I�x$�W�����;�C��!E����<��|'��*��N1�d��@Z^�^2a��M�m��E����F%4�/g��L�����������_�9	�7����}��N���(�0i�59��ߠ��H^óor�Cv7���ޯXĜv�_L�_kԊ��n۪���l9`�6n������[P/�(��?��iN^�W�+7!ρ��E�
�o2<����=�g K{����u�4���&�I{t��3g�����x˜a�q5.�%xs�^�OR�Q߆��j@ ~j���<�,}Bt0	m�j�1����z-��R�EH����	�<���֟�}�7@�����j�� ��9�E(��n��lA5�:,i�$~�&�\�+]�!F#a�,gA�c���)�&�H�3)�"EͰda�J&Yf&E�h���ۺ��P�7��Z���\��0�^2��>ؗ�|���5t2��}i/C���`��n{B��6K������Zݎ�w6�?�Ӟ�ܽ�E�P����W���_i��'d�Sc�@`�&9�2*�0F�d��)�6B���$�VF���;j�JM~Q̽�����Ns5.�{_��X<���ˡi/w��� H&}<�i8���"ol\��nJI��=0|N��o�;X~���'O��^G^�*ݩ�YϏoX.]���G�膛O,Y����C�;�'c��X��9�?��`$�)$ �?�d�`��e�|�����V��}sG�9���B��u������������"X�F3�j	�.��դ ���y��7ހ�����!���ǽ:a���g��{B�[_xeZ�[�wW=Ut�(v�l�1i�[��[�XNA�o�w�r��]?H�_>�l��/�X͹v �׃��E��)�Ǎz ��վ��x����{7�"Ŋ	�.�'l�^�|G���o�����׿iq��9jf���B�ĸ�SwJ�&��zK�x�G��{�o\�S_��>�Ȁ3�Zr�o4:&\�y$�_(1 ��8XeX.�
b�$�O1��Ua�C�!ؙ�|��c_�|���'�p��W5bYC1Y_�a2yN���v��O�nA��E�������#��4-��yu0���4*���lm���)萯��#p��x�U�yl�u�����$[�mL���p�(�=����o���sJ��B�Șv�����ȠT�kH��Ƽ�U�O�o�_Mk��p#��!R �GpO�@�Ɋۉ���gmڋ_}�������?�/Y?����#Y+����啽w�Sr��_�~�d�%�z����!==j�&�� k����E�1�}-F��͸�{�۱6��!���Yn��d����"�t穱#�~�8;�c|h8[u��-^�bŒ���
{6��77���^[K"޿���+_#3ӳ ���C=3*c5K�S�O��EĴ��t9aE+�N�ZE������֞$'���>��o��<�}�V��$��t�^��`�薔����|�ȞI�b�v��`/�>��^�����;_<2��e��,Y5�Hȫ�*W�U�ͮ��ԇ!�v�0�z�&o���
�i�]+�t>�cjk�7�y��y[T�e��\�x�2z��w��Q���E�Q���k_���5?Y�o�'!&�c���r�CX^�_�[�y�es;J�Z��d���ê�v�G.MU׹3Zo�[3���o������f,����{�N����^ö[����=�l�+�0F~�\������bOl�1�g���+����7O��f��!�BϺ�'M�S�$Uvq3{���Rd�P�G����)���	��i�u��3/T�תWq�_��6?:%gm}��6�v���s�!�C_�Cb:�Y��t0R�������[�r��b��Nu<ٹ��-�e��!�`O�փ��im�Z��ܥoK���"M1�?q2�O��t�҅K׬]6i�Ϳ'�̘\3�ea��O��颍���;|��;��~R�ַms(<l�~ü	�p4V�G��/�������])��{��1˳�G�h��Q6'z�(�b�:���7r5f�qJ	��թ�-\Y[�mWş^$���C�k^�S�R٫aǤ�/���|�0����?�!d9mz���!F��X���0��
�3e?��2��՘L��+#�.�/���8���M��X��ƑA7�\50�I�YBc<���Y��C��B6'�{���D[�ܑ�d��ړ��?v�7��/�_�gx��Ƿ^9I��Ρ/�{K}�|���?P_޿�/6i�P?7�:"��C���������O=���E�8z7{���mNR�jݺU�׭[}�_w��q�����W?����׶��_�_��ᮘg�|�c�H�	��x�=�mc<:���'�A,,��S��nI!�r�1�Y���<$������Z�^���lZ�1J=�~a��(�����⩠�E��;JM(f��i��1�IR[d�^9-�o`��E�FƄX�[�mȆm���H��Yc��PN���{��Z�n��[���=���������;x��=6���kk�*�F~:�������)��~q��}E��V��k��	�U�lU�1H��ii_j�5I���:j��Y�gU�;����ʝR?G"�"ɓ����x�Z�1oθW�._]�nơ�S�f�^�!a���.����4c��`��[��<|�gϜ��׀���(d]�7Hρ�w��u�n�r�'�L���#X=\�Gٺ��N��W��y|m���I>ޮN�P�����aVzN=���f���;�$�����܆Mh��6��I_gCa��������ґZr%4n���j��=���W���؞]x_l|��Y?oߕ���f�\���MB2ʋ�{.$�>Z��C	�2�B2�OJ��OT,	%(�1�/��:~�r�	���H!��$�����8'W˿��I��\�}��]^,�=&�g;���Owf�e�dŠH����p�,��Y�L�*��f��l2�ox�qQ;��Y'��j�?�^����Ff@�iM�2?������9���4HB�Nr'%�f�KzI}�JwC?K�!ɘhji�2�2���B��
���<�t2[�i�k,7wu3��  DL�.��4������F���B��4�̧��|6[�k�o���wo��?l���N��a��C��/�
�A����?א��-�]�A��A�f�b��GVd�C��/p  ���y��=M>F��	�k���9�af ��F�r��k�i�}=�灶�/(B��F,+��P��g)2����m�f=Lc�H�d4�`#��"l�Z�k����Wq�Zzw�ؤ�oj���@2�����3������&&���Յ���->�=�>����fE��nuquq�quu��z� W�*唻�IOw��?Mz<�\<�!C�LF���͎��e�R�._�.�N������������=�=�c����Qe���O� �7����9A�+�m(~t�`5�NƃOႪ���蔔-N����H�U� ��x@&�'Z���W��5~��=8e��A���s�M(�Rb:{[�C&i#�ѳ�Y�I�E�32�"��� �HV� �AV�e����Syr'�̾����z��3M�)x��<>����3�'�kՐ���!�����8�~�N/;%���?olU<��鐁B�k8i��ۨ@�2�HC��]Z	�W�L�Mq6�r_���^�~Cԏ4^��]'�fV;q�C��R�u��E�5ލ�'�d�H[��tsel;Ȯ�z�\���&�� ����� E:�w�����~�'��LVS.j����L�V�+�e�v_�t�.�\��ֹM~��x�!<����Cx�!<����Cx�!<��� \��?����O@�®��f"r�u��p��	b����4�3���,�B�������[�����C��u�z��^wE=��"̌pw̔��1����:A� �N�ڙS]B��az]Fm�9z݀�����E����.���^wE�����*/�RPi�����6y�-�����</�8̖T�n�-*���^�������y������#�l9�%S�*l��y��[Y���[niqva��OFvI�mxiIi\i鴑y���%�����1���/-��*a���ʲ興\h�^^QZU���_Z>%/�$�2bF�ܼ��eeɅ9y%y�b4�K�(��cE^�mr^Q�N���{���4xζi�5f���/��׭��̅����<;7�8�|��4�%�)-����B(z���\SʳK*�r�l�� <�A{a��R[v�,[��N��K��,9�4�YY��";'������@�HӴ�c�PIP' �kˮ�(�)̆�@�9U�y%�ٕ����"�qGNQ�e��W� �u��畕��V��	2�� X���<�C�a`����\�Ɍ�ʂҪJ`��P���/�T	d�*�?'�V�'���(s�#��QZn��;@�B`U��Ԝ9 [�]��NL4�������U�%0a��[j�(�UTM���S�[4�Kr�rJKr��&S&<ʞ\:=OH�y�`��	JJ+�Z+�JY�h�l� ��<]k�8yv39KK�/�mť�y�V9�,/?&
טj��8{�_\�[�_�-��\*@4;7WH������r૪(�\L��WQ8�D�1�hVYA�=4;�T�~*ZΤy\����"'-����4QK�f�
��:�T���I��
�Ln������QZ�[aj\�A|n�[_�ABm`=:/��8�*�bzia#cy3+a�ز��`�eO.��4��r�dW�
�+�b^Is��tM�k�����<�i��e+J�����ʶ���ѱ,;gZ��bIic�����l*Z�b^Q>gjH�-15%Ӗ���9*6=���aKKO��o�̀��0ۨ��!�#2m�#=6%s�-5��2�6,)%>̖������aKM�%OKNJ����A�#�R��`\Jj�-9ixR&�LCuRI	�����AC�66.)9)st�-1)3��L������̤A#�c�mi#��R3�F<�MIJIL�Y�'�@hPj�����C2�`P&4��2�c��Ǧ�����6�%����|pƐ��d[\RfFfzB�pޗkgpJ�p��)�I�)��%6.9A�D��4<�;<vpBF�$��.N�:���	)	��a����AI�zLJO�)z��Aɂ�A�)	�����2$AL�¿A�3!~
���d��g6�2*)#!�����YHLOv�=a�q�/E�ۈ���Ћ���O�M������w%���+�侭/n-<�P���0�Z \WkU�gXYb��"\���[r�~y� ��H���� 
V�P룔��b��6X\��{�E0�j��2��U4��|A96Ĳ�B2�����-�
Z�g�[q��U����Ғ��2ة
���
���|?��@V��.ԗS툡��)�x.�Z�̈́A2]�f�rT���T�l�#�A���"�Cm2���8�S	�u%��C٨�Ak*����y� l(��V��˃k��8z�P<Ԧ���
z�@�l�2E��A�ӷ��e�g2�-�~6_
�f�g-�d*��p�U%J)����0�TЌ.�����;F;�6��/Z5�*u鹄��_��3Թz���?��µ\��[.�y0&� ^�A���3�i�,��d!m��'%:��Ѝ�F�ۄ?�,��-4W
�u�_��p�S�Y�s6Ԝy���L�Oa���g��᷶ߐ�PעM<�V-Z�m�����,M�+Ԛ<V�] ���rM���t��Ӽ��4k�&�*���e���f�?MT�[�Px�&K��i�J�E��-~�{H�N�A���x/j���ZAN^$,�-ւM��R����P���|0��XP�O��6X�㎍<6����ւ��|�&��2��0K�೉�\!A����R<u���3��k)8�T4��>P "D���b��,��~y3�Ը�:s��{:lݴ~+`t�/��(g��R6AY[�B]�ͭ��R;4�q[��ѕ-��I�Bſk�j��D�0�i�\��a��51z�zZg?.ң��B9b�\�q��i�X����l�X*"C��cQ��|w��WCE����R���<�&d��-5�1n;|MӆɳŞ�bG��/׼��ڼ�,�o���vx3M��X��Y����W(ֲ#�q�+����h�r��:������E�WP���
N��J��1E��߅+gr��l�=��:�h���ߔ�9��6�la�q��4���^�c�n�"1��W�z������:Z*=ӱnZ�"yz��kf�B�\1>��bP��-G���]7��۴���b��,�}��U�zpXb:<-|��xNV��5�w���e�Ț�8���Ͽ�b
D���k��c��_�M��p��J�"�����JP3��k�BDOǞݴ�+�gE�9H�>�9�2��� O�-��%B�-��/"�/K5Y_#����ߨ�!(A̓�R��ϓ
w�h����)�s��d$��?Q/�+���Ab5��:���FZ�t���hh�m����)@��M?c�g�TS�n?��k!I̩�)�nF��QHA��F��R`T�X;|�E�4ڛfm�U�����p�K�C����B���b�DQOi�3Q�4V�S�4G�⎷��k����2kܦ�&K��@���� �]�E�� ��>S��3LH�.~X����g���y��J��K�����3g��lB�Lh������,(o��B�X��T1C�xƵ�����3��*�����8��b�X���J���:����|	BSɢw�1�'5�h��$d��V������N�$d�}fM�}*V讹�
��7I�Y Vǃ�t�d�ݺ�m�*��~��k1A���h�B�X��u�G8y�Î#t�Lm䬹~��������c������s�Ѩ�ߦ�Ů��r�yG��x�k�s;g�MY�s���b�s&�E���oq�~M�Z|����3�s����qJ�r���ב}h�[;9g��"O�r��ƬD�?J3��iӞ���E��^��W��Jђ��_f�l��V� m����X&�{m��^�g&\�*�/o���T\��T�[6p��[�/�.Cڙ�Ph���:�r�8�5�k@{/���՛��S�F-�P��)N�����W�s������q������������D�Pv��~����ed3Զ�-P�<���P�AvA�E��"������K�U�&'��:9�7�P?G�A�<��0�˖"ʖ�w�~�]��e�.��c�C���_q!��}[�[^A�R�	\2���ׄ���H�OL�D���ٓQdά�"4`Jy�4�V�]jC㊲+K�˄&��Z���H�
�6��вN��,z CR�p�1L�d���&Nu��>�1,�c��HI��"��a�(�V<E�WN����`
X�HR����|�B�(T�:� p-���o5�9���L���'�\���8W�7=�i���6�5�=���_̈�,�k[�	CBfz����:͖�P���H��,�Л�cH�ı�9��$�[W��l��L�m�ϭ��^���F<�cT��>	���i������g�����΅'��H;�F��?��>��ˠO���Ɩ]��0�54�ʴO�Kï�!�h��b#��"!��l!訥�BK�X9�� � ���5�9����]�FL�JZ��$�t$��&1$�$�t�E&�\2����d.y����g�I����#��r��O>&_�o�Mr�ܣ���B=�/���igI{�~4��)4����h>-��t&}�>IW�ut#�J��]t/=H��,�Hߥ�O�u�-�E��zF���2/֚�X(cQ����P��F�ql2+`%����/a���l{��`��~v�e'�9�6�®���׬����2Ub�I�J���R��Q
�zH�R��(%K�R�4Aʕ�Je�ti��LZ#m��H5�Ni�t@���I���%�}�c�K��t[�'#Y�-���+�����r��K�'��C�9S#O���"�\�)?.?)������vy��W>(�O�g�����u�[��|G�W�bP\/��bSB�0%J�P╡J�2R���m���
�����T��H�=ˁq}�E�[� �kx��>W�U����	
ɀk�'�;���uq��p�}&<]'�-�&��~�x��x>�=�^��F�U�s{G�B��1�Qr,�u��h���tj�\Y�.��Y}�y� �_q=z��j�x�}"`8'�� '
<��Z#^,Zb�-�
�%Z��-�~BPNx��Y�c�[E��$	<J�d
���!�0�2�c��7�c �OGr�?���L`�}�����q�=*�Yg��!��I;��Yk�}^��Z�%��h��O7����d����aM���h�u`\+�V����&a�Tu;ט�'`G��|��������w���j�ǫ���qM�"��,||�I�����C�!�%�^	5�k��v,jQ�v,�h�߬}.����o?�|�jx�������p�jz�����6�Q�ml��LՋϥ��hOlN����:�/q�����Ũ�4�����	��-ڟ�o��*����٫�>վ��U�8nxpNAk'��a�r������������]U����?P����焉voa����'��5+('�!�#�>�Rx���$ֆw�ӆ�Y�e���S���e�V ��J>J����L�9���m��Cęi�C`o�#�*��Ql$YcEZ�^@A�]�� K*�t�tA�G,���8� 4Ӓhٍf[�@��K�K��K'�N�K�0������ۿ��l����+=[��U�Z�<��i�Sd�]�{-�|&}���-�DKS.c�L}��؞`�ؓl1���[��H�=�(���� ����P(����D�3�����Z
���
d����ӗ�,�����O�u�-����zB���/Қ�H(	#Q�@��P�FF�qd2) %���&���<M6��ଲN'��Qr�!o�+���|M���.Q)�&j��h[D;�pڃF��H�i:͢h.�J��t:�>A��5t�Bk�N�����=M/�K�}�1��~Co���CLf��|�?k�:�H֋�cqlKa�l���Y+g3���d+�:��me��.��d��	v�]d�٧�:���bwX�D$��*yI�%�*�IQRi�/�Ҥ��8i�T �H��li��DZ%=-m���vH����!�tR:'�-]��I�K_Ku��]I��l��r+��$w���r�#'��r��%O�s�r�<]�+?!/����-r��S�#�k�c�i��|I~_�X�R�F�)ߖ�)H��+mb<��x�$�`�^d��޲��H=����\zp{^Ƿ�����IC����	�g��P#��-�,}C�2���?�F�:����H.u什t�G'�	�^�\m��B�-	r$�N>-��=�2ioqʤ������O�J�2�.�����1�����(����(Q�QNx��1g:�G'�$����d��J���H^��� 8���EK����K&�S�x��:��҇��Z�c�� �m�v��}�h�ώ�Gp�%��)���o��Y�S�Y�O
|������B�������?J`���w%��
����F?
|O���$�-p`\+�VQ�HCo �CK������xޒe�;�*)�׹G���#m)��0��q�R>�.��O�9��}�Jx�B�	��*�T�9h�"�H;-�|�vKP�{�M�x��4����Rx�$�c�c�1���8��>)��g�J<c�q�ؗ�=���N���I��郿�l� ��A�[&���oS~��I?�����j�:(�6R�;�ԏ�3t�@��9���9����&���ɥ=_Y�
���:!,V�Ǣ~]��ۼ����ZE����I�K��S���d�py��#��<#] �v���[�]����K]$���D�z�Į���� �'x�#��/�{h1�^²\?�d+_Ar��K|���ܚ3)�}Τp�׹��R��-� #�x5Z��� Qt6���hp��ly����-�|�Ix�(췸��SO'�ĩ	�Z,e��[C�_�^��2�)��9�h6r�q��P�<{É��^�3E>�+���YXbQ�%2�� �	B��t�|�S��|&���w����Xc��Ȃ�ė����3�$�H?G���IƐI$��r2�<N�$+�:��l%��.����3���"y�|H>%�ɷ��C�)�㟮ԋ��6J�h�C�x:��ёt�Lh	��������O�M�9�����!z�������
�F?�_�:��KUƘ�YY+֖��,��`�,�%�d�β��˦�26��[�ְl�a;�v�ղc�4��.�����K���n�{�d�"yH����^�,EJ��~R�4DJ�2�1�$)_*�ʥ���ғ�
i��Q�*m�vI{���a�tV�(�+}(}*]���nIw�z���U��[�69T���>� 9^*��#�q�d�@.�+���y��J~Z�$?'�w���C�Q��|N~[�"_�?�����仲�0ŤX�VJ[%H騄+=�h%FIT��t%K���*S�2e:dqO(˔5�e�R��T�(�Z�rZ��\R�W>V�T�Qn*��{d������oho�l�4�2�3��RX�S6�2�x����TQ���/�z�}�Vo+�\o�;7՛�r�����x֩�S}�3�=�4��h5*damDݹOk1�$��i�3�*�x�F9K��X���/��j���7�p�y������������O�Ug�C�����_��j�O�>�I��S���]�X�|��&=8��cm��ޫ������y�ΉS��m����G���-�_"��t���O�%����9������Ǧ_�^��<�tjѢh����|������+��m���$)���v'
Yb�w�t¦�w��6��;�=D���s�$��H��9��N#�9�x�=���hڄ���JB�Q-���(�FgP):���������+�7�=�����AwпP5����fd�2ڊ������ڇ[� �������Wq/<����@�6�	��rc��01�h~S�~�~��/�b�|�|+�O͟a���1���I�\.�o�O4"�i�5��{>�P&+J�R��V(K�U���&�9e��[ٯR�*'�s�������4w��UW|���}����h��"�E��a�#�HiL�4@����Ɣ"J)�)bĔF�#bD��)��2�a�R��0�aJSJSJ�""��=�^^&��d~{9w���{���{wO�j]]]��rD6dO�.������A�Py��%g�9r�\ ɳ�r��P^*�`L^�X#�����&y��]�)����G���)��|N�(_	�p�0��pJ8-����
��Od,��(DLG� ��E�e�x�,�Q�X��ClDlFlC��
����#���G'h�����Kx��XDB�G4�I����7�3��p#8Í��Ep���ɏLuG��"����#����*�ZD-�рhD4!�#�#{�x qqq�i�\��e�5Ɣ "��z�>=L����S���Bd+9J�R�!������AA;Q�"V(�e����Gl@lBlAlG`��Q�Q�I�#���)�rN���
c�� _� 	X���A:�x�^��(L�"��P�P�E�?S�G��E�V�j��uP�;@��6؁�.ʇ����pN�Y���;@ݩ�;u�j����=U|;���TQs�x7aj�:N�7{=5��Sg��9u>�Gݩ�UԜZI���Եj�Z�6��3u�6#v#Po*�ME���7��� ZUԜz��G�i�;{e����4ԝ���Pw�NC�iC��Z����h�Z�V����j��Bm��B[���j���m��Eۮ���h����#�q�vF;�]Ԯ�Ln�)z�������0}�>V�O���B}�^����"}��R_�W���:}��Yߦ��w����C�Q��~Z?���/�Wɐ�p�T���۸�h1���8c�1��7�3�Rc���Xl,7*�*c�Qk�F��d4�����q�8i����q���0=�����c�7�C͑f��m昹f�Yd�2���Bs���\e�1k���s����n�4���̏�#�q�y�<g^4�X��b�eY)V��n��X�0k�5�oM��Bk�Ub�Y�"k���ZmU[�:k����f�vYX��C�Q�u�:k��.YWmɖm�v�T���۾�h��ۙ�8{�=�η��3�R{���^l/�+�*{�]k��v��d7ۻ����}�>i�ح���}�	:�p<�������w9C��N��͘���E �{�^��A�u�{�^{U��A�u�{�^��A�u�{�^��ك@�u�{�^�8�y��9z��^좥���.z�k�)n����s��0w�;��Nt��Bw�[▹�"w���]�V���:w������pw����C�Q��{�=�w/�W=ɓ=�s�T�^ODo�~o�7��ez�	�$/ߛ���J���o��ܫ����^�W�5x�^������z���1���z��޵�`r$�H���'�J���>�5��ģ���������s-��謂xM�e&�ӑk;���r:�~���C߿bύ�[���$/���ʉη�r�����z߆�y��x��t��Du�����v���;�F��~GR��;\r�k�=��>��w��J��-��������sGҌD��U����ڨ�t�]=�mܗ_���qk�=�۾D����R�_���F�6���>y��'�'Ҕ_�����.�:^�ѳ��m���s7��l�:�k�]~[��<�Ȓ(�O!y��oD��2	{�Du�l`���WW@< ��m���XGF�D�[�����<�3�o|=�5��왮m%yk�<�<�,�v�It�m�-񌥓�m%=�J�}I�7�6��<O�=O�l��9�Z�&.Oq����(OY\����G�;�������D�K��&���|�3��1N�Lʓ�L�P�!�'DW%��ўx�x�&��v5(V�{�?kj6�Oў3���T�S��g�Y�_;���+(OE�������/6L���N������y�TN:]�@���_�/�'�Q >�x*�OM��D�j�m�D��r_Z'�l�5^��������7�H鎞{���b=�؇1S{r��M|4���ˈ�_M|���r���x3��G�L|2�b�����c��!ލx�_����c-{P&��(I�)">�䃉��=�i�g�B����Zt7��Q�+&^ܮ�������ǚ8�-&^L�A�� �Ӄ��Ac=����i��$]��'�1�X�;VֲA��mg����Yl���}�<��o���K�i�?�?ɼR�w|ޕ_�T�M�%��\i*�F�)R�4�Ϡ��%�9�g����xy���^x-P�W%%'%��I]���/$-IZ������o�Ƅ����P%3�|�y�1TZ��
U���&Z-xGyKi���w�F�H�[h�`��g�$oR{�=x3�g����kY��Uz[���(:��e�GYҮ��W�"AG�U�3�s���+,&$�� �B� �ا��t> �s>1
G �wh<B�����8&���*>���J���T�;���^ �f�w	���ւ8�O+I���Z'��ӈ�����z�/!�Z��gzgk�̂�? ���i+�A[V�u��o�=R|'���F���b��U�*��ZV�X#kb��G{�v�c'YkE?�̮� �p�{�;�����|�G�,��sx./�E|����B�����^���|�����ž��\������c_��`"�]r	�[�`"�P��KF���a�������!& ěU>b
ra=�x{� #D���X���O�n?��ٶ�hb��ㅔ.򥅷��y{{Y,���#��ρ��Eq�S(�>+|ќ�"?�bq�2�SF�?�����xOκ�	�XSyxbO�3��	��y8S�ͣ��<�ͣ����Gq��).4��B� ݏt�},�+���X+$�:y�46|���sYfQI�6nzq�d6���x>����,�d���s�Μ=��������z�==Z��՜Di�F+؍�.N��x�
Ka�χ`C�H66k:3VR.�����bO�X�>=�����X���qe�|�W�:)�WI�Tt[���(R�u��:�r��Z&�l��M;���;�a�0I����hd���o1�����c]����!E��̣=����cen�=@?7$�6�qM@D��e��!�#0���	�&|����d�3�����|~ ���	�~/�K�+x^�7�-x�Q>S���U�����$P��dp��BW�
�}�"�8���\�3ڮ�r��O���Md��x��o�w�{0��<x~?��O���<�����Uxބ{�]�s��o�?�O��!��V�C7�_���s���#�E��؂��X`zp���v�g)��E,M�Y�90	� �@)�A9,�E���JXUP5Pu�z�f�rAiQ�*��s�.���\�THk�_���	�A�A;�&&���~c��2�z"W:ك�؆g�-���FL�y�}:��μGgn��JEQ4"^�=��"��(� �Ox�M˕p����(�=���%��7<o�Cu�?��kD�}��b�y]
endstream
endobj
20 0 obj
<<
/Filter /FlateDecode
/Length 448
>>
stream
H�\�݊�0�_e.�������@.�C�>�c+Y�F6�s����#�C�8HG�q�v�0.T��S���0D���t�1��4��RT���n�*����⯇p�h���Wڼ-�AO��t�_���p��?�1��}�?�Շ�jj�9]����wWOU�=��?.����w��c�$�c�m�z�p����v���|��7�ӹ�b>��u�u^�P/P-�&/G�J@�AI�=�T0�0P0�pP0@( �
j� �*��U0�*pU�[�`���%& t���Z�fiÛ��)QV� QHox�t˛�w<��<�Q<�1�l8��s@+8���*hKhT���Z4��4Ҿ�(�� �@@�7��y0W�`�DAY�#e8�:�[�J���`0�t�u@r�<"e�aYg�s�{�i����[�n���0O����_ t��
endstream
endobj
25 0 obj
<<
/Filter /FlateDecode
/Length 14941
/Length1 35396
/Type /Stream
>>
stream
x��}xTյ��g�s&�B!�W	B��~���$$�2�LH �ę�����R�R�)E�Q���R����-Zk�U���"ZK-Er���뜙L��������b���~����k���r�q�X ���M+�x����5�����O�N�Hc�6�M�K��~��?��!T/�^67��i1�0v���aY��ݽ�1���Uջg�H�c�h��U+�\�
�؀�hsku����F�_�X_�Z�42�Վ½��nu��}�[�X�v�xݞ(�����S�����ϸ��~@M}Ӫ_<���Sp��:_�������|��ֻW5�ժ�~�����<~f�mq�/�\Ϯ��	����m,�����;G�R�9��ȍ���<�o�o��7�r6t�P������֪��sԛ}@����9��D)���,K'֥ q,[Rc\����<�4ƴ�ڏp�l]��X����h����~�҂o�|BrYIu����+����Q�?\�����i��Y�}��?dc�ݬK���h����e|(�]ǮgO� [˪�&v���g>�,�
�g:��e[ٝl/;̚q���q=�汕lۅtz-d��x�2�PF��aװ�]�vX%zo�})�[��#�c;Y	ڏeA� �������c�'YJ������rCy/���-P��}|<�e���6`�b��m`$CV�C
���M�b�/�r��$CrYHa�DH6�^Nr��t't��$Վ��"ӝ��`i�C
�cј�Mhw p#R��,2���ȶ#T�S$�sp�@����L17���]*�O���Co�t�I/��Bf)5��=�07ɹ��au������d%��d�R�l}X���7��Ǻ?<�B�-�&�~�b �� ]��9�� K�K}Iy/����,1h������$�MTڃ�6���>>{�|���(2Mf_�F��\���Г�h��/Iò��vIjt����Y��y�7�jdf��x�g@o���g�iX9���`U��7�xv�F6� �2��u~����KX������'AI����~���0�J*�\VN+v�e������0z���� Y�38�	)zc���氙lz���l� p;��̣���g�A���]�>�}��P��P�x:���.�o�=Ю��O7_�}�@>�s�����a����m��=�b�B��1�3v/�z�_��}�/��;����_�y|"_�˔a�A�woB�%�^��Q_��O��S�<z�3�k���Ř�'��!ׯ�����������xC��g�������f\�fK~�0�^�ȝ�����~�u�ݝ��JXS�0Q��hƲB�n�f+q/��e�� ���Z��+1����,�eS�J�l��jY�9��`n�1O��`�ð�*X�jE����U���m�t������[��g�d	(i���}?���B�Nȭ4c���n+F����t^VH@�P�X�*=�ȮB�X�#� �G>b?q��Z[t���{z��}l���-���;�&x��(9 :�C4���0�CN^;a��K��T�&y�J{�n�~<�^�Kw"Or�V����oi�c�F�;!����6(E�9FopJ�F�Hy�b��N��t��;]%Vn#�䗁n�>(��(e!�B�l��j�3�占8��bem��l�TD%%�-��r�/� ֕��0ڭ�jߋ1���=܁�ܟD�� ��~�M3h�A�J6�e��R&dt�/���^��}�a�H��-D�eG!��O�/&'������f?�о��$�a���pv�F��%]�8~��A[S0��Ak _,?¶`�^`�ZAc��т�n�����3��Om�>����l4�i�����_5�e1R_P6K�/l��qѼ�GO�ο���<�h�=�����eG;連.𩽨ă}�X	���W���G�lܕ���ao՘�X�M�a��Y��3x`0��K��{�.�y4՛�n���ߩ�7`  >7�w�A�)u��lDYw��EMwV�'����:�ff�n �
i "��*�e���<�����Zo������3�C
�%K�R(��"#��X�Q�B���֬E�R�X
��4�"b*Jr�J/(ES離�KET�1G�i_��#}�L2.���d��Pv���5�R�쑱���"�[�S�Ɋ�4�t��u[�f�:st�<����=�p��/�|��֚�1�UYnG�����Z.ll�hU�A� XU,�����7��G^h��f�s͹�uep�N\����zk���_h�p���r� �L}�2��/�k�wɫ��7<�(Ү���2~�,�i�6��6�|���Qt�)}�\��t��~f��]~��uRO�7��L7'�YX- y�bQ��7��V���W�sb����X�o��\���jh8��Ea��A����l;�g��v�;��cq��^�w��qfd��{p�K�݀�D�ƾ�K��)�A�(� u�����qM��i��q�!�_���a�H��(Cd�E�@>�%�4+m)�x5ۈ�D�{������щ�8#?�ώq������pO\�w��;�O�sYAD]n8��`<�%vK��D�E��5=V��sVk�jP#��mGW���~�ڈ���9H��}eе=U�Z�~�QVB�������T��<�Y7�]����`	#5�8��a��6N���g�s��a���`~��9��-d�Y��=;��T>�^�����E��)B�{S_�?���"h�v��	�c��tB%�kE&%�u�	-��Nuv��?t�	�/ӟ�Oe��Zp�#v˅��v y�8��9m+i�1�%>���i*g����S�ů�!�V[9��� 9����`���ǚ���]Fm�W~�`�?Q��}��c��=�8��?��tր�紒�_���yU�$�/�z�ͥ�C*�����|����и��_J��$���2�VCt�tyPj-<�N�w�5ħ~	� W�u,_��LB�%��|,]�%���h��7�Sl�0@�Ys4���	��M��Έn��{'�G��}n�.#O]��[���v#�m���F��.A<�f/��&�d)j{�U����۱��v��nXg��
��O�F�Ql2����������g4⬵�����p�Y�V�uL�-Y��N\G�T�G$������Xp�	J�p�c�Sf��<+?|e"���6�3A"��8%�ǉ�+����b0�C���D�� >G�:�]��
���4%[�c=��-8�e�������F�?����z¿A�A�m�� P�c@a8x�ޮ/� ܍ �����$}�+�Κ�S��'RP����P:D��_�s���7a_AKAvt�؁Fз$ռ�O�o ^f���z���Di(v�2�1�e��� DJ���y��*9����d�f��`�Ѱ�4�~Q�.�Y3Og��h$��.<��=����D~�(�#�v��w������<H���
9ؿ+��<
���*B^g�.��|�W�OgO @�?�7��ǐ�\���?��*a��2?�^���z��iu�W��/w�)w�L8�J?|2|�|(� �t�]�ς��+��)�����v���D$��q�~��#��|���{[��� tّy��j�w���I�9�۾���������X��{��VNt�kX/���ː����g����6�TN�/	�\�~<�����6�o��ދ�j}G�>�Ň8y(�'v]��C�v>q�Y��]8^ݰ��$��� 99�?g�Ӑ�|����iN�r�Z�*|���C����Kx�Rk1��i�W���US��[5�/�n}.z���1�7�� )��([I�<�NÑ����>���HӐ��IF�v*$�XI��g�R$��d�\�vZ w��Vr���t����E|s�Y_����Sc���ߡM�}��>�Y"e����u6����}~��5U(�e��*����s*\/,�74�í+��:�JvZ�:�T�����Ej�A5���o�<14cVI���3�y6��%y(+�@Vޡ��yT'=���_������]qw��pW�w�PvDY��t�O=%�|J<q^��8��t��S����P�x�E<�%�-��]����]����!S��y'm�y��Nb����������ڃŃ��=?K��,{�՟��ݦ�i���M<�s���)8|=;���I��s��I����,m�r��,�����΋�bk��Tђ$�o�-���)6�b�7N۴V�{O�vo��gc�vO��'�N���w��Oiw�b���O���;nO��X,��VoO���Y��������E�l����>K������#n�*nlk=�2q=(^�%֠��,�:I�B�*�Xi��h
t�����L�o��2E#j�
_�h�Jk0E}�b��)Q�N��M����lu�r�7˞���TQ�>5���Q�����7NxLQe�JS�׊%���#]��-2��	ba�X0��� QT$����6���\S��9��8Q��s��1�$N��(J�D�)�f{��1�#
M1�3�j3[DAW1㼘~^L[+��j�kE^W15I�Ċ��Ĕx1yR�6��&:�I�b�SL�]��"Əsj㻋���qN1.[;&I;V�sc���QI��Yb��mT�� �F$iY1�#���aIى��<1,Id�(3Y͈׆vC�(���jƐ�ZF��8�0���,����n������u����YbPg1p�H���������I��H靠�d�~�QZ�)r�(ѷW�ַ�H�%�}ФO�� z����E��h�g�x�gW���GTg�G��!y��&%��D"�%��ncE�Xѕ'k]ϋ.Y">.K�?/�P�%:�Vh�׊X��V�N �)Y�Κ�,��Eʣ��YDY: ��)a��kњ#�#<���E�g�=T�E��&���,X��p�m��!��?l��ܧ����v��gx[Į@�@�HQl�j��87,�[-b+��iԍD]�:I�V�(���&�!N�z�-^�P��&�ee�րS��h� ��=8==���,OE��<����#~Sp}����R����0Z�f����uP��{��`o�3�[�V��-�vW��я�	�����γy��������`G�je�򼺄�z�8�,R�W�������'`�[�6�9�څ�,ƪ��{�����`���c��bojo)�q~��b���)����c�ˇ9n�Πw��p����j��Fۍ���zf�Q��QZ���aǎ��⎟>~zx��~����ը�B@���'��{�K�.����b��z�h85��b��F���K�qv�KY�9hH�q�k}K"�y��׃��^Ȏ������jrL*��)����㻏���11�`�6lҩ�c(��Ł���(<;�#N��#N����)�n��|qvi��ѽ��J�2Y�*��;�u�Î�c~��ULlw�t1L��9g��J�����&qG�����'⾨��w�Į��я�_��QOF�\��:S^��uPúq�t�׋���/�������G��?�4!�uʦ�C���垯�)�4�����;?�n��a/���n�F��=���ѣr�9��PMU��<��ݳ��lub��t��:�&�N���5�`c��=��,9��Ξ>{:��Wg�����.��e%v����S�n	�#�ƌUSg�4[��x,��Q�m�6ͽ/w��!|O������ٱ��{h�+/a�q8s����z�j	�gMlBM�?�N�$��,QɊOt���)�����>%���2�,��R���.#�9�3zTx�� �a?�>s�w�Y���Qw��^['�U��qz�����I�7����ȑ]H��E�k-VS�O����n��f�6u��a�E�{�HM��%2#36�W���ܝ�p�V�鸏�ĝ!�g;_5^��j��^�-�od���/�K�	ңC-�>�����O��?x��h��G�c��)�F�*�����[�]����ٕ��<�*^۴����2+��O'�
���a�N(�k�t��&������͝��'=�K4��艮�t0}��iܱS��))v<TK:�����R��Ǔy�����'��/��E��<����-.��+��[��ɓG���Jn��~������Ϳ~ޫ7�|��"��9�㸅���m*�}=�f����nFL�&�YW6�T���q���t�؅IǤ1����
3��c���7%��]Px�y�����%֟8�����Z1�4�^'���EcQ|�h���V�!�]86~��c<�'$N�rJI㷘�S�J+?5��~��)����W�6�xǒ����8Yw�?��^Ӎ�t���?):�K�H4ғȚ-k�;3�����qı�)L��]��v٪U��y������g>3?�<�=!���w���Ϳ ��Ǟ�ԛ�vӳbDtK5�w�c:E'2g7HvZ.#}�X���,����j�6��yUo�~��Ӓ���C]9)0J��ș�V��zA]r`Im�ޤ���w��~�=����:�&GE+���ɩ�1j�3��ʻݝ�:�&��ߨ5�w��%G;��r�)�c�:RF��"�p���H�/-9%��[�9�%�����!.���������tg���)=6�밄a�2�{��ION���o��n�y�u�U�y��ش1à�ѣ�@��9WTz�v���������ݿ�f�Y��ٻ������:9�F�?�$K$��|�/~ѿ?gc'L?nRJ��]v���0#��+����":����f�԰I&�u�M�{β��$̐ms�l�����G�M����'���y����gf�x�]E=��`���^]�tV����@S5�k��T�r��`�9θ�%�1�{���SY����e'��*t��%
m���0M����b��@���ͱ�zqu�������������Xx-bYhM�ݰ��By���ƌ����M�E�=E��+!.M�ʻZ��ϊ�/�SƘ��f�K�5��`5�fٽ��T����o���I�s>�<��|��q>%y�-p�;���d��?ǟS�E������E�p���W�
\�+p���W�
\�+p���W�
����+p.��'�ǆ���,�?n9�Ý�W�3[y����Ո���d�u֕���Q,�}��;Y���w��>{��ǲQL��F��h�r;ϙ˙n��e�.W#�Kr��y��9Ct�X��{v��&8�󝺦��|,�q>6�׸�_����5�*ݕ5|�HW�jWnmS���u�g�
�2]9uu�R�*�*���^OfL�w�{^����ݰ�p��^Wm����������ջkBm���l_�ϕ�������WV�ȱVY/���j�O���5������	ÆyP��93�k�Wy�}����oӰ���k��6x��2k��Vy�i�[�$�
���z]��:���L�w� 3&��3w�,�a����'&�װ��ȵ`���w{��n�r���#������6@�E��ߋ����M^O�����C{�&��ݰ�Ո�@_e�mX�Q���l�T�'�]U�oDs٠���,M���JR�A��r��Z7ƃ���M�&�Oumt<HR��2_u�J�<%�8�{�>Os���xj!Xmes��xh�!�TU�쑜��m��57���Z{ ��o�d�h/��p�{Ij��@MF�r�a>�+��<�u-X���0�dd���l��@+k|�w��P��o��^����W��r���I�X:��IJ��|�Z)G`BLL9�ܕ�^���"b l�&LC�*����fV�+P�P�^[k`F�n'��v�w����K��jZ��vc�L������Ւ~��S[]+�]��CD�In�N�/�|5׹�4���]�@l,�[�X������@$ {��	tɲ8��0w]�D�~!^�(�ņ�ծ�v���^��7j+3�L97�%��y-V����+%�S�ء
W�\�)�6̎��V��ڌy�B��Ն�jªq���ܕu^Ya��&����q@���^/���=�f�H����~%Œ�r3�[�ʦ���v�I��j��Z�^
����C��V�������Z25#�5����UV<�|~Ni����URZ<� /?ϕ�S��������s�]hQ�ST��U<͕S��5��(/Õ_QR�_V�*.u�.),�GYA��¹yE�]��WT\�*,�]P�����&U�_&���/�:�9���2\�
ʋ$�i ��*�)-/�:�0��U2����,4�@���hZ)Fɟ�!@hjqɂ҂�3�3Щ���Ҝ���9��2$����EM2�%h�����e3r
]��e��9�e[���Eų������r�!JNna��D�Z�S0;Õ�3;gz~Y� ��-N�:d���E��9������2=��O-���=4QH�N-.*˟3h2#��� 9�7�8#� ��S^\Zfe~AY~�+���L�0�����D)�\�SN^�ͯ�#Yv�u���m���S�e����º�WUy��mۋ�r��J-��AVk9���,\����g�,�y,׶�䖜a�_�>`�؍,��Y�HW����dem�V:��z����u�­�/�u���~A�6�F-����6�����(�׮��b��Uu�@�ґ�7Ј��v��nu&���~F��6 
��E'�U5M��&�R"����2]1l*�!�^����-e5�]l�b�f�ထ�U����M ���^2���ր�����E�Xi�V�z�{�2��!��f��B[7�,��.�%}�4 7��{�pW�;��GYבNQ�f�U��ه�����GT���H6��P�P����ǩ�zK�&[R�&�:��L�c�_���h�������O�f����z%�Z�4���}W��4QVH�{�3/�1vHO���x~d]���ZΡ���s%�������Lz9ץF�4�F.���-��P��9�����E�Z[�.�wӬ֓V���;�6^�d%D����ٮE��꼶\Ki��Gѩ�Zox4k�-�� �|�a�o�ׇ5�T���%��d��5��D\�_n��"i���(���u�lZ�VJ����̹i-�k���B�-�e�U��z��D5!�T�1[v<(�c��SH���,;�#��D�4�0J3��ƍ�$h"[�/m����<B�����Y3Q�t��l��<D���z*��(D���*-n�I��#��4���n[����92�r#/�"��z�h��Zm?���:�9��ưE7u��6�V�>����PM����1���#����JX/$j
����:�K�f����ǵ6�hu�۽��|��� ��i�bO�@�o��@�����xI��E2�홪�퐭Yڰ<��2���e�}=]���ٖmV���$��v��\_���a��i���Zy4�{�����S7���m�#�.��Q,}5�����$��r�"���^�(w�@x��u��X���~�*S���07�ѥ8�<'��먗K�a�{����W���K�շ�*	�-3�n:�"^��y���J��C�S.�/�����C��)�f����L%�{_���z��
��^Bc2&k��ٺ`�bn��p����x����!O�k���K���bIw).k��(2R_)��WR���?�fv��%	��Њ�D]8��=�Sl$�^�Ԟ1k_���������f�*�5�d��aM�*�q�Y��8Ÿ+g�O�R�|ё�^t^� ��G��C5�>�V�|�%�bz�˦Q
,i/@���{y7�@K��g4F>�PI�,%ڳQZ�k��N������{���d4j�W�^�vd?ɋ�i9��Fm�U��l6�JA�]��DO�A����0��lNsHG���9ҝ,��k	ڕ�>sHf��"�a�-Y�k&,���Z��e��r�B�Tn�� 	�<y�_�:�J-Ί�Y��6*��.->\�:���H��:]$9J�inr@?D7d;Ӊ���%�rH�4B.�I-J}�[�F��Tҗ�7�y��C)��$!j�g�R�a:ɗO�*��e�c>��K,{, Y�ں�hZvo�Da�v���rf�`�|ۦrHw�V��M
krl<5Bgm�_d����\��]�����U�uYX�h�ζ9�aa�y�k�gq������P���;,Z����`�S��aYX�N��]��ת�c�k���߹#�Ƕ�42��`m�62���tj[ߡ][�埭=����]j�
�����-�E���F�ѯ��t+��k���#��T۶�[��zjy�и�d�v������Mт-p	m^n��xBl���e%���D��l���k:���NU�6!Y�M�~��Ff��jI�2�̴��Y�|֦�뻰���f}���1�:X��Ǟq�{59f��v4|�7қ�/��2�E1%�ߘ˘�>7�ufB��qe��#�)ې�_�1�;��WoP�`Bݠ���k�kȿ������ȟp�d����S�22n<ba���W��2�]cr�v�}���i��,��wW��U��ul�R�w9+�s�\lQ���JSI� �o+�����a��4�DF�G�8��Q,��l����E�����B�"����٨�YeSI�X��$�F8�~y�r�c(�C���)L���d�r�%g4K`�� L�(6	�.H'�3�k���a�%�7[�����]$�ji�'��}o�����+�Z�}��	���,�G>�%Gkɩ!�$�ߖ:RoVo�U�7���[Ȇ�]�_��)[�s���(_��G0��=JQ�d���7�����<.Y<
//�F湲=�;\rC��&�u]�$!�%�Z+.C��p奠�eY"#	oT�CGI�m]!���W��Z_��~�����芡tQ��de�2X��Q&)���H)W*K�j�N�+���[����J��]٥�U(��'�g�_+/)o(�(TN)�*_(_)�"�D�H=�K���%Ɖ)"O�%b�X$*E�hMb�X'n��U���>qPO����q\�+>���KqN���ƨqj��[MQ���(u���NS�R�B�F����FuV��X������ԝ�u���zD=�S_�*[}O=�~��QϪ�5����EKҒ��`m�6F���j3�"�\[�-Ѫ�:ͯ��n�n���6k-�vm��W;�ҞԞ�~��������Q;�}�}�}�]�=J�����KO�3�,}�>E��g�%�<}�^���z��F_�߮oԷ�[��n}�~P?�?�?��������?�?�O�_��tӡ:bq�DGoG�c�#�1�1����(t�:*�8<�e�F�
���g���R��B���E&�]�� ��
�I��@��z�z�P���pF�_���3I֚��>�|]pk+��_�qE����E>��l�B�{�|X�W�PKp�!� �j`��W����>�����PI���ӭ���T���cp~*\�Q���Δt�r�;h�"���U�5�pq�\CW��nne��V�cJZ�u�٭����;�Z�h�d�����(�:x?���v�˒�󩤜��r�YT�Xb~<�Y�����R�<���q�[啄����.k[�KYպ�t�Z�|���fm�=������A�N"��k�A%��X�q)��#>��g�����?�ޡ�<�	a~�-��,�C4��.�k	�fN���� ���<�xs"Z.6���|�4��0~ ��k.�sM���%��	�?���3��/x��F��e1��a��yp����r� x7�����s�+�Si���՗į�~~�@+���(,&�#*y�������oA���7�6�M�n*�ʟ�%wt�9Ĺ��Q>"�<��?Z�cw�A�t��rFz����H��G�Z�[�,��/���!򿠖�}�k�,�s:07�I��7X,k�V���b*�.5F+�kJ����W�?�6�I'HW?��Z�����c���H�`�Kk���גg�$K��$Z/τ�?+�P�by�����Aʮ�4��x�(4b�Q��r]Mq��Y
bLi�7Ҙ�H72X��dLb+���=W2N���3����d߷#�W.�l�et�cn��M��%U��J�G��P��o�tI[d�}|-�o7������!V���7�YoK��2i
R�ޡ+{g��\uI�%��c������f�*w�;�����Og������(J��$(=���d(Y�8e����TJ�y�"�R�Q�&e��N�]٨lQ�*;���>�rXyZyNyAyE9���|�|��V�T�)�PE�����H�D�%&�l1M�RQ!��L4��q�� ���mb��#��G�qT/�����=qR|"Έ���T]5�.j���P���1�$5W�����Bu�Z�֩~u,�V�.u�ڢnWw�{��!�I����K��;��S���W�MѢ�X-A멹�4-C���iS�<m�V���i�Z�֠5ik�u���Fm��Uۡ���i�����s��+�q�]��#���vN3uU����D�����3�Q�=[���z�~��ї��
��f}�~�~��Mߩ�����G���1�E�5�m�=����~F?��w0��0]I�d� �`�p��$G�c���Q�X�X�v�9��U��:�rlv�8���{h���hw˼�ų�kCye�(C�+�܉z�r��R�
�G]�oȾV^�a���
��?R�s�,�S ?�;�o��Q�g�ԟ�c鈔�a�+�_��T
ɉ_î��,�H�U��2",k��w𷅌�V9J�*[�W�J��T�G(�b*є2M�nP���V�j=�'i�GO��+q����E�ܗ�'��Ϗ���&\��&<�p.�%��Qe4U�Jyq8A���Z��ƚ�Ӯ��I�\�-����j8�(��
�p�㣴s�㴗�W9dT�������Q�b��CF�i�.�!b��}�:UFz�ޢƅ�o%��Gպp��D��2���Z.?���r!��|L�^&W����/��I֪a�c����s5D��Y�	*9+�#JJ��a�ۖ�U��)�r��oS��iQO/����B�a�&m&V����N��Z�Ԓ&�Z�-w菑�I
=ɮK��L!��4��Y[��U�n�Ց���9a��}��x検G~R�3?��V�*�w��p�*��+�~m��y�zQx������m�u�%�K��J鲤}b]�Q��tpF�.��oP���"�_GdB��Iq�F]�C8S�}
�e
�����O��y��It�'��P>�����!�{:�cvB����%'��>�>��ه��T.W��bc%Fr˟Ԧ�t��[1G��p��G��d�1W�L3��<�y�-�r������P�HM�s��1(y�Z�$<��1������Y��,ii��,���"�BI����B����2�xx���G�|����r��/&
��!R�ʛDM��W�L���G}8�K�Dm��}���s��uy�����ˉO�pQ>����W_B��#��j EP�)���"�f��VW�l���8�F��>�8����(C}Mz�D72��<���D���A<���x6��y)���p_��
~��o�����6��������?ʏ��k�m�����t�5f!�~+�#<���;o�hSsQ�ŵ�1ߡ�%�K$��Qy,"�4"�f���s�5�\}�<Q�)]d�H�P�P���|.��~~�?��H��r��@������3�	�+�8��N{��D貝�9��C#'ص /�:�o��]�L�dNlEl1�:�x���#��rF��Fs�wbc䋛�8��s��=��u�:��?����/�K6��o,����Y��32��3�q�'�a��l�X-�e����>��]l�c�c#�ulrlb�[��刉[X�s�s/�9�9b��_8��΃�GX�y��8kv��|��t���[-��NOW=W�º�odlR%R���h����uH�#mD���"���H���#=���H��'m�?�qrV��N� +N��(S�;�;O���w;d��v@�}��0dyr��w��#v;Ϲ�����!���L�%�M���?J������p��u��oj�]ʿ)9���+�>��LO�z���g���|�o�Lz�/��in�4g��_&˧T���%�^[�|옿=k���{֘E��ѳ�
z�XI��"��=m��|z�����v����W��Ss�]�$��xzN!0=���'�����@V��
zYIO +�	dE�I'sd�p���NFW�^6�SW��M��mp��چ�&6nVR竪c�/��zjY�_��a���~fi�C�%u���w肰v��V�����z�ٷ��ZW��~�'|�z�Kc�S��η��|B��I�4��B~�׈8u��m�y�4c�Qh���<c�q�QiT5�2��h0��
c�q�q�q�q�q���h1�;�]�c���8�<������S�W�3F���F#�Ht�FO#�`6R��۫�֙��؃����g�g�\���F�QnT��%��h4��U��:�Vc����l�gl5�;���^c�q�y�y�������0��8#�`Fo�e�!�VX��Q0S�Q���.�YQk��C~�:�k�G"��ɒԟ�o?m>���2c�q�q�Qe����Ҹ޸ɸŸø��d|���q���ƃ�@�a��ο:?v���w���p���Π���k�C�)>8K�K�d��)�L��s
��NB�@�����Q�g<�m<<%\s�jQͣT�F�'Y.}*��+v~\H[������K��U���ö����]���ϥ�Y�����L�
endstream
endobj
28 0 obj
<<
/Filter /FlateDecode
/Length 281
>>
stream
H�\��j� �_e����n�B`IYȡ4�$:�
��1��}�	[���ϙ��3��}i���>�z���:�0�4�3�J���)���n[<έT���\���p�f�`�N�Sz��w��VkpF��uǐ起o��������W~;�_��f����F�b{���Bu
���V��?h$ɆQ�z�󬎆_�ɋd�G��('z"�D"
��g"JV�%�
]r��{Y�WR=N�J��)YY�F�ǖ�����saT�{Ҍ�t���Zc�*�_ Dg�
endstream
endobj
29 0 obj
<<
/Filter /FlateDecode
/Length 622
>>
stream
H��VMo�0��W�< *E}E��h��mv���r���a�$gR�m�!pL��#�)�Y�
N�v�
(���[��(������Ga<����N��G8Y?ē�(����w�&�B~/�'��6*k����{ 4 ���]����3h�;���6_�S�h��ҟ�gc��BϘn���O�8��s☴B+�{RX�����nB��*�L���b���G�4 �������Lb��5�G��E�i�gf����E
�.¥䵢dr�ٺ����n]��5gZr��� *���c)��	1�X ��V��\|JY���[�﬊1'P����٥R�͆� �J�D�k�+�m��iX�x��.}�3����0l.mQ9?��UziM+p����x簱�潂MD�,�}�=���OA�K��ս4D���bd�Jǯ��0>vsź��N�p�v��\Ytm��[(4蔊�ʵ�):1�0��;�w:]�)K�m[VlWZz���i�$4P�����D
t���8��"�ja���v��\d_fv约�]�v ��/&f�����G��W������`+�9ԉ�f�����N��M=z����G�7l�!0d�����%��t�c�J'�pF���? ���
endstream
endobj
30 0 obj
<<
/Filter /FlateDecode
/Length 553
>>
stream
H���MO�0���>#1��	U��r����j�� D��?��#`��l�)�M������q*����'&��{f<��k��M�W�;F�l���͐;���-OW9����Y�{��J6���/���7f���n�w����>4/s$����7I�q�dO�!���Y2W�wf�z3�,��S�U�)�΄���٩S�i����{��{t�Z�̞��.41Dp4��N$�}>� ���6�P~�ݏM��SKXs�T�<5u��5(]��r|\��1��2G����G��խ�j��X��1z.�F��7qCf�2i�N��`JD&�Ⴉ�-�^V���׫�l��֝Fq��Yy�������v{�"���@��	�j[8~�^B���Uu�>�S+�u�.O��b&G�Ns�ZUԗل5���"�.05����U�[A��`�M��H]�w]qG��<,��6mm���f�ʓ6��!ݘ�'1��`��Q��LeY<=�A�1��hGQ1���Ӿ9d�8T��ťn���R���~���/���/�'� /��
endstream
endobj
31 0 obj
<<
/Filter /FlateDecode
/Length 496
>>
stream
H��VMk�0��W�<��OŁRh��� �2vtc����&�uq�:�Fz+���8O�O�����^�<H����N�X���_,^�'�iŷ�P�J�5�,c5X_!��m/T��ϻ�){Q��d|C9���ȣ�!v�Y��n�쾋�=xg	��"%͢��p�`p.�����3�������Y�fy���`�C����f�2��@�M>��W���]���4hS��֚�k0�*�|�����Đ�0�!��9�ntE@XaMl���|�� �A�ǽ�ϗE�����.¦$tv�)���^�D�-T�J��� E�^zȒ@	W�Pu@�����e��p���Q=�l��(m�<7E��TyӜ����_(�o`d)�8�6�#��������P����:O}�0խ>i7-����D]����.�Lפ=�8g���t\6B�đ$*�"��D7�@�r��$�D��b�}��=f�5n�x>�#~YB�F+���+�	VI�~ �܍
endstream
endobj
32 0 obj
<<
/Filter /FlateDecode
/Length 503
>>
stream
H��W=o�0��+�+�t�/�T!%Q�n�آL�ڪj����aCM�4M�!�a��w��A(M�|p��@��jŗ�(�����W��7F�s�6�?K~P�'�kė�tP�[X#��(����Mp��(�i|����7�G��U<�M�v��C����I����i.Z�vK�C�H���X)3�a�@�R��?�i�ec4H�g�G����I>�T�����r�>'�3F�2H��e��T,�T��D�lrBU�lF�BN����|;��㉫��>_ȗXc�<�*�4"pOc����G��ǳVVP�EKK��"�!ciɮ�]�Ɨ�3���4�xi��ش�w���ې��D
�.������'r�x�*��q�scғ�@'�褷�UjR�׾q�K��m^Mk��~�aS��r"�;���i�)�C��L0(V_�T}5["���-���e ���T�tr:�\��:�f0�]Z/�tJͰ�m��M�駌v'���w:Y\}(~ �A��
endstream
endobj
33 0 obj
<<
/Filter /FlateDecode
/Length 519
>>
stream
H��VMK�0��W�,&�)Ȃ.z�&�&�q���$�%Y;��FJw��}y��e��^�N�S�n �.S���A��y'�@�׫�Wv"�h1�ȁr,>�!z/�A�L�uH���kx7F��v�
 �fz���=�%��%.-��z������2J 5Ѓp��xk���x����i�V�[Hf��M2u���x�-K��1q��/�U?�[&h�u��h���T���]F_)��R�K�kt⒣��ʸ��\���RՀrdMt��ܲ:P���>+��4i���Y�ou�V
9ϫ��bK9�f~�L�rpr�7�-ch\ ��O��ɉ@�'Т���EY�Ӈ�B��8ĳ��@g�㽄J�Bf��M��t���Z�.��ƕ��R=���w��x�2�YL��-��&,&���=��2�3:�_��x�?���z`��5{4���v�PPk
p�Si;���),`����Z檙ag��)#���l~a����<��`�ת�6$�������_D{�v!�u�BRt^�-4|0 �\��
endstream
endobj
34 0 obj
<<
/Filter /FlateDecode
/Length 475
>>
stream
H���MK1���9f�Y��-��M؛xT���L��fu�M�TJ�YH�y23o�8���C�|�:��-�Â4�r/x\��gv�6C�4��9,H0�k--���zxc��}|o^��J�6\�w?��!�-aU����C���"q��EԴ~���(�-�NP%gSL�1~[M��^�X����)�u�L����Vsl��<1¨~���G�b�:�b�)2#B��s���a�#x�QG'����x8R�����z�P�YؗQ4�8qS,>�� Q4��v l�Ӷ��2.�E.�@�W�Q>�Ѷ��{��U��9B�n
�'��s��G`�VOөmZ�j]Z�d�F����Ӳ`�5�L��uA�`�*���aw)[G�:[w�(��U���J�������F	��F֛���p_]ld�F��\��|U����z-6{�]jv��P��L�Uv�=Z���S��).�e���	0 ]Б�
endstream
endobj
35 0 obj
<<
/Filter /FlateDecode
/Length 467
>>
stream
H����j�0��y
�5�b;�BS��n���N�m�����a�[{�[�uGi����gK,ȟ���m�Z���>�+(��}4o�S3�~ ����>��F%�BiŸm��`�\X	��op�|���|�]��#��^j��2%3�<�����c���Y�d�^��~}���������ݭ��8A51����,JU!�&0�:I�
�FN`r=��8WB��ʑa+�� ��F�O�i���l�\���B���-L�'FzH�D�5��L��0ٲ�Q$��j����(vQ9FN�F�dk�@c~{��Zfrc$����\��u��C����A��䝟�z��lY%�V;)ϩd~g6%̐������_�-i���a֢~ц�;V�d�b�G�K�O�Z��ߌQ���ďuU�u��q��>t�5��L!���� �uP��)^� s����p��]� G���A�
0 W��e
endstream
endobj
36 0 obj
<<
/Filter /FlateDecode
/Length 489
>>
stream
H��V=O�0��+<#�t�؎#������1!Bt��?p��6�qpҀ�ԗ�z��㝍�Q��4�PP���7�"Į���xC�-�j��l��w��]Z�y޻��k '9���(���׫���rr��1~���T�e�*Pvf�%����i�g�x�5��	�|JHCCy�̺�E��iD��G_������?�O��8��zg��&��F��n�
u,�UN#'��f��G4*��0Q���	��"��D}%"�Yf���/E�E^wnV�U�-�dWA=�0s:�����DIK�ݠ��k�-M|�TX��,a䏕��-�~�X��cխ?{�2�S��*��]��������(ܜ�,�H�CRA����ꐭ^'���%5K!g~�uüf!.>�=(7*���Ʒ��;_kƗC�&>�tW�>����r�5ƫ=K��9���Q����A����t�=��Qc��1-����<�h���o ��1
endstream
endobj
3 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 4 0 R
/C2_0 13 0 R
/C2_1 21 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents [29 0 R 30 0 R 31 0 R 32 0 R 33 0 R 34 0 R 35 0 R 36 0 R]
/Parent 2 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [3 0 R]
/Count 1
>>
endobj
40 0 obj
<<
/Count 1
/First 37 0 R
/Last 37 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/Outlines 40 0 R
>>
endobj
39 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227162545Z)
>>
endobj
8 0 obj
<<
/Type /ObjStm
/N 19
/First 141
/Filter /FlateDecode
/Length 2623
>>
stream
x��Zko���_1m�� v]�F�4�������*dQ�h���=��]r��R��h�9��ݙ�y���cM3��lB(&��c1YJ�!��ǡ5�)��*r��!θ`J��xoj���䍏ȳ5>#���h�35[|��f3�b��~��׳�?n/����K�����z��|z:����\�mn?�'�/ֿ,��������J;{�L�>�{�߭���/o^�.7�Y���\ܼ^�.ݘ��l�r�EOB���������כ/��1g'�Yy�1��h�\_�Z|X]�߮�W�k����i�bu��9��|���4�����?�Jˣ�	���jq�eN7����_�����ŕ>|�=�}{�Y\��?���Zb������O�Bz����8s��٬�濺Q�P�Yy��[�ر�p�>ݡ�7��^��cx���>�t�ק�HP�%ء�~���̙5g�b���`�A2�(	trdM0!fA��$2�W�^r0���X�H`�a
h�����Y59��ɤ�r�Ho����K0	Ԭ(zЋ�<���Mvm��6�VX�g�KB�5OhW��&P4��c��3O�7���@]��c��<�[�^����'�U��B.&X��yA�rM�7Z��w1�9H.s�y��ǱL?_���Lh�OD0WD������g��m����,��q��vl��q?������� 8��L��K���t�������-<���N�Fy�������g�z!�Ad��@��'�$��e !KG� H6�d����$!A��t$I�.�)D�=Ǽ�ް�Dξ�s��8�P(<�9�t��	�-���*'.��)I���͙��+SA�B�g�my�,�
|�)��b�+W��U��L)UۯXp6��a4	k��H��e��|���H�vb
��`-�y2�p��lY���C+RB��b�K�Қ%�vh�,��IT����͹������B��<b�g+-��X�,>'�ʞ�I�,i
$5�#V��y�E�w@_�gP��YB��oAۥ�5��DG�ᶉ�f�C���J,�B�	��1� ��e955h��n���� �@����$V $�Y/���J�"�I�ƊI�2����fO��H��{h����:�Y�P�)d�3����)��,4���4ǐz9�=�h%O0���zAE��� ��zsH��PT�X�C|#�}X��wЍ�*vZE�&!45��Jmf��zI�eqU�X����/� ���|��G���&#H�2F��1�c���4C�U+ԃ�K��5���>[���Xh����\Q{�/�O9��}���(6k�m5�rQmQ�.�bωv���.ζ���Q�!0*b�|;L��ؼ�'�O�?�~׭� ��c�F>�(ʽ���d��w��� ���c�#�s�_�����N"ne��!�� .��_�%���iw����\�ں�N$�"�A�4C,_h������kl���R�av�R��
wI6�j-��9��˲Z�L��0g�P�CVkςMX����u�ֶ�y��i��^��!��<�v�Л���q'���ʉ�'�UҀ�f��R���q��� �w�B��~�
��Q
���I0����t]��=�� �n[NE�T��A%�T����|W�"�
�oJ][%�Ot�)H��@v1���j���g��B�y l���N�Юj��)���0���?���M��>�_�iwj��s!|���"����`��N0�0�.u�t�\���N���)5n���k�~��ϹC�ݑ���DU�` RxB�����ajJ�_r�@�c����<�*�� ��1�Z	d�2���-��m�er6Y�Da �ݼ�0����!�V澋Χh�㵈wU,�C��Zj����m-������v��l��
�Xy�� �E2|�����Ǿ�nx~FD1Dj��N�q�ā���N��1��%�i�%?�c��G<!N�L��#���@SFJ��}�Q�8���"T9��6��p(z<��"�>�<%��`�=� }a����<��:}�O����kj�!�v��s�:�ou�s>Be�,�;E8�{	�����R�_N��z�*��^��ߠs�C�|~�ۯ�̛��G߂����zÒw&�E�_�߯/x#9�o$O^���{����+\PA�n�Й�uf�yvBGy�S[
�����ry�I�NR��~�I��$Re�1Q��U�1�$I��$Rd)1���e�xm�Re�1Q��~*�A�H<,Q����ps�uy4�ui�(I$ɩĨE%.�H������h91�"e���I��$�����T��D�$�Tb����*q��	D�<TRI�H��TJL"e&�xx�Re�1	,�Hܒwa�4fuw	��+w��g�E�/~���]To��]�/~�������7o^~����Ƚk����{W������]�ݬ�]�?�k����9�d����s�Х�_j;����󍃷��8�H� �w�=D�E����$���	����`�����qL8�&	�'���A8_~��Q��ǐS3�f�v��0g2�x�ڼC���_j�?:Z�������8 �t6�~q�鋶��쿍m�
endstream
endobj
41 0 obj
<<
/Size 42
/Root 1 0 R
/Info 39 0 R
/ID [<51888BEFF55B2B4F9AE414499E1C2ADE> <E4FE5AC74F77E08363A97A3C4A92EC12>]
/Type /XRef
/W [1 2 2]
/Filter /FlateDecode
/Index [0 42]
/Length 146
>>
stream
x�%�;
�`�����$j-x�6�^Cl�A<�� "H�v^@�!v�q�m>�vY Ue��rC�; B����H���3�X��峎h��hY:�"m[|<�D"�"��ϋL�<z�㛜f�%��f�������oa����#
endstream
endobj
startxref
50463
%%EOF
