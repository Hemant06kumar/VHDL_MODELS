%PDF-1.7
%����
10 0 obj
<<
/Filter /FlateDecode
/Length 23
>>
stream
H�:��� �����pn@� 3
endstream
endobj
11 0 obj
<<
/Filter /FlateDecode
/Length 2818
/Subtype /CIDFontType0C
>>
stream
H�|TyPY���+fh������JTtaF]AG�@���G9�
����@ @ 9"�C� � �*�
�Q�x �%�:�ʪ�[N�v�-���g��j�������������ǁ�@gy�����u��D&��և�SU��rGq��+*\	z%��hM������
���ޯ��K�h�i?W�KĮ�U���z�q��ɒ��Db�R���ek��4%�����ˁ���ى[��͉�^�fooo'nv�ʩEEhJq���'M�ɳe�D�X����̤��
J.V�幎��ġ$
J,Q���T"[L���r��R�E�Dy%sT����+J"�X-*J*q�%����������,SI�r�X�a�ވHM���D��.;(-���\h-@�(��CP�p��!(��ul��e�2�dàph���wY��w3��E+�xB>���� V�3�Ղ��Km���9,z\���e�B��
�i�w��dj����G��P�p�N�8�`��,
M�1��w����O�;s�E�:/]ſ��m��5R^us��G�\�)e���/��'u��!u5�r�ᘾ���������X��\T��S ����'�ȓ02������,hmm8݃=�����L�p�'��s`���ʺ���� �oᯐyZ ~C�ךf��pja�Lh؅3u|dF�����x����@�@<s���
9�7p����c���&��Ҁ�����l"Lu֪Ny1>$p��ƅ�OGG��<�t�cu@�_9y �u���B;���~å{�5�Q��8�Ÿ�� x=��g �qt���1�.�/��Z?��ÐL
�	�0��ɩ�m5�dK_���4V���s�<��^r��c��ӆگ�b���Α%����U��}rzb�)pŞ�ݍ%&���g\<��������V=�ߚ�J/����7{`̖�ń��> ��+�e�}4�;G;�� ������y�|� G%���M;ѐGj,��o06��ư�B��H)?��L�	_��ޓ'��S]��FҢ�S�{�?2^)�݉-��~�P_k܄-|��y�	$WF���3m�M}lpCa?��?;�J����(S���c�08Q�U�%�L�g�|�v���"�Y?� �v��&�Ͳ����5;��8�bxL!�0+A��#k������l?6OVU�0�4��n�38�Ms���R�PZT���5M�Hp+���C����Yxx�~�L-�+*.)Ĕ6uKc}MsQ{�l�XuM�m��sI�I��d���y9�q��?���wt��Q�o*�	J�ۏ5�G�4i�9����1��u��l�mo�c����Q��Y.�.z�p��(�5ȷWo���zI���X��[���Fsq=i)H�$㢐��h2(:=h'F���'�	���{+ao��h�D��j�󿂢�N7^A3*y)U��1�~�F�
x��ڸCژU0b�UJ+�pf#d8�_L��m�2�$����Èl����Z%@���IT�H-H�L�%�������i�0�My�pf@�.��*I$��V��`I���T������{t�7:*�p�tD~h/��� �3wZf~ �`�z���r��`���"�#🛆�Fp�������?�z���֕@e�y�j����'[���G���_):�ޏ"o�TC�!� y��,M7K��?���Ky$��h�:#'����2�\h��T�K��Q�Z-(,<����O|�pq�,~���_[0��>��Z��Ѵ�56�4����-�S��/c ���ɳ�׍<����f37;��%������E��r2B|�����aҺ��~C=��N�G{J.������.���u��	�g�XM���I���;�o��>�z���t�c���UYe�
UVv���F��P|��7���K8A_�c��Fi�W���D,��*B��j�73 ~��ۖ��0SY�����]�����<_U�.��	�x��Jx��d<�1�𾲲@=��lp����"�@�z;/�:��%���z]��Ѯ��>��3P���t��,���1�G�-����4�7 �1�5�.���j�,�	�X]M9T������$�����?׎w����I����[v_Z�uă��I�cI��M�q�z�>������Ká������|�ȑ�����������s�i[`SYm ��!������������ƃ��vp�b/OPE>�j�o�t�s_aiofO^��yq�g�G�}|��x�����X�@�^�c��������cP��=������������}t�rrj�������������}�JIB]pn�����<�cʔ������v�;���0�\��q�I�FrĄ��|[uJk0h8n�c�q�{�������ar�����Q���������)���֦ǔ����������!��6��A�5�!��o�N��f�)�(������ԯ���Ȓ��Jr����ykyjwlwnP�y�������\r���Z��n^pcoh�cY��M�q�O�W�������������	�p��`�q|��v�1���3�V��r�I�Iră��evL`�
oG0��~�������_r�~�T�D�����z�~�|�~�vxht_wrlwz���{s�s������������4��9�ޤ��Ĕ��� 
�&�s|��I����%���������F�_	��
��w�n �U-
endstream
endobj
12 0 obj
<<
/Filter /FlateDecode
/Length 293
>>
stream
H�\��j�0 ��<Źl/J�j]A��M�b?��49���!��~1�t�����Ir¯�s���a'Ѡ�^iiq�+:�fqR	wW���5���f����'V�?}pvv��EN�����n�f�Y������$���kk�����C-}\���k�2�V���t1I�M+жz@VD~�PT~����S*�z��ڐ��(J�rSrJRJ:��Hy�O�t�I)%�H�B:�*�KP�*����̩g��N$ꙟ�%�ٮ�_���~�������)���5�_�}�W� vf�

endstream
endobj
17 0 obj
<<
/Filter /FlateDecode
/Length 22053
/Length1 48848
/Type /Stream
>>
stream
x��	\TG�7\u���+Mw��� �!܉Q@@QD�h��,�a�h�$\�[��8>&q�8�!jԨI��$&�$c��>�0��1�c������РYf��������έ[˩�թS��	%�8�d�JN�S���k�ُ��#��}XYN��Ax�;"}lf����x�L���#2�%L^�v)!�~��SӰb!�E��[�S�p��|�*&���Ϊr]�h���IB���%I�|FH�a��=#k daޭ3��P���t�_���gp���@!�u��<�w+,���bO�@�g���Ą�NHb!��Jr�;w���e�*�)����I�L9����*�܋�CX����+��c�:�.�7t���Ե��9��w$�H���{��>�_�H�#��x�;��J�.��{߯p(G%�����G�	���͜�2�
�{t-Q��Wٌ� ��>"�,��eI��J���}�����Hq��j�@�J�W�����X�=R�y�"�4�!]�`�Nw��d'ɦ�h�B
�r�l"�Q[��J�YH��u$[�҉�a�J�x�����ۤ�#2��h��̕$��#\GN��J�%t	�ڃ���ypB�}� �'��rt���t&9�uOn�Tp�G�h�/Xܣo%�	C�[t(��l�������L?���{%�<��9�^����x�F!�6�}���{�7CO��y`������	B�BPY�TV�շ,#�w)�
_��d�uq����A����f?j.�Ш嬨��d]�TFY��.�\)4�\�`o�s�V�O��w+��-'�q ��u�!�5�L��F��%Y&<g9�Q�Hg/�Q*<�>��Ep��Om���!���1��d�B�j+�#`�-��?������	�s}�����&+!4y4^ߤ!N�h}@萏1b}�C��X�;o9-������GXtv�����Z���Z23B�9BwQ�-v�y�����sm�j��Qrz����<@y	0����G��y�� >ͽs5y���Z��R�����X5���(�3�}-��;�9̂E����f#�?Jt�z���a*y� ��حߑP��{r ��f����|����o�x��t3�A�9h=}p�~��I{J���й� �7�.�Q���L��_�0��N̉�������'�L@��3�a��4tC�x�>����������3����ަ�Ak*�7�1o݄H���#�p��\A?�dp1b�81b%����%w �����$lU�H[�����;X��;����� ��G�o�G�?�-<b����"�>X/��>x�dX���Em#��r�o�m�$�*����O<m��T2�L����0*D+'!؇��;�j+�s���L#O��&��S8��퀷��-$��\�GZ����|g���NB��)
Iv
��b��h�rɠᕎ�)�$ҥ����{CđT��=J�s����Ԁz��B���/0?c磾 T���ǥ��.	���K�ęd�P�8!F�0���ƌ�\�鏕�Fyl&��/@�ǃ(�F&���z5h{�3�^p��V����y�x�v��[�*B�<5��������3�,����7��x[���0��!���x�8�ih�
�D_W�qڟ�������<���Ftx���;��E=��t�X�0y��}�H!v@!��k�:f�Oy��#~I�����AFR7N�� ��+>D�!�@�QB_#�($+bЧ(I�,�2��>�����G$w�� �`$����Sh��Q�Dc��.`2v��b),r�� ��): �?�U�|@_5[�y@�F@�;�e��=���PRL�"��OrH%l�,�8���2���'�e� Xi�Ç�_A~��&���nIr_�l��T�⾆�j��8���'/�D��m8���b���<���݆�,Om%�A{)����Y��K���X/��@�����LAM���@$���J4�\B[,�=�00���A��af6J,Z�Ї�m�t$"�C4�<Jc�jї�8�y[G�o8��X�>�Ya�6L�z�Ρc�Y�B����)����^�م�x�*oY�y�fVW0ƛQyK ��\��}����Z�R�mISi���1�(z6����P6u��j0<e�Ȅ��᱅��̳�y\(���8�y����&<��-|m�O�=��Kr+@F�k��Nn��u��kx��н�qe�J��x�)��{�{Lc`G�Z-W������;ڝ��	,��h���j{�=>��r�i���R-@��IZ`k>1�@�yE���/�Kg�8/����S/�'e�	Y~��-���B�
�����w@�f��*diw\7��/p~�(���Qw0z��&�'��!�1~�_M+j;�[�t�CF!���]=�n��{�[����}���a8M�1�i;�ȃ'��,�_�}�&�T��?���Hjż��GT�,�c@<Z�;����ab����A��ax�1Q�Q�h�VW�G�^h����8�^Lp:�L}__�%Y�Qb|��f�w�w,��c3��hI���J� M}��������A��1h��z�v�h<G��K���TK�+�sh����-ȷ�߶�q�}ۚ���(��(�}�}�,<���Ž`�ව줽�	�8�3gn�;<���ǝ�0��O�? Z�GZ�'�1c�&���٭��' ����; ��gvs��d��[�[�i&y�ȾcM�{�ȥ���+�Haď�́���dɆ�;�"Qd�h_ �Qq�ʦD�k����-�m��m�SxQ����P#��[���q�Y�� �$��U�%#��Y+�mT(��t�v����P��!Y�����T��\�HO!����9��x�>���^���/�z:�9t�wݻ��)Ѓ_�9.�m��P����H���z9����>ջ�' n]d­ۚ�?�ơ��TU�'zW9#�E���3~�?~��|�e�B��!��]�c�)D�޸9��G"?3"w���t��m�y8
b:/Vd,FPHÍf.��AN����	#:�ӈ�V�译�m��������.��n���8�2��c���n��f����KМ�ەbp3��y��8g��;�c�����ƭ�n	����Af	�"��@�2 pW�[�bܚڐv��A��(!�տ'|d,��]� ��A�G�-�0c1nrO ��q�=���Z<G�ng����mnb�QBQ@��l0��c0�#jѐk ��z;@z\h�gO��O�����Io������nBKnD�HD�xйF��Z�L?���y��耛a&���b&� q'�&��� :�ߣ�îpv�՟F⳪a�^���9��l�	!g5�I{Хt)ό�[9�O����Q-���,~�A��vO]ێ��⦐�?3�_S���V�<��17و�,�%���<��� z8?�I�dG���o<�k���a�P~Z��3��Oq���'��x!f�����>�GO$���/v|"/,�G�J4�x~�'���t4���x�!�6��)�~�?��e�|��i��O����[@��<���٤�`�������x����8��˫xB.�W�w�t��4��^d�ޟ�N��oM��ߔ���7� ��7��"2w�NJ�f�C؁`���C�p�{���3[\��]��?���>䟱|*���u1NA��98!��߄a5&jx��2b&����Ŋ8�]� 2�1�])F��K��^r�1���@$H�9�-%�n�����q�w���U�ݱW��߿��U����.�-[OJ���%%��)�xJ4!��S�m��WB�<c�=e,J)J9ʃ((sQ�AO����|��/�,_�B7�7�_������>�yd��X<z�9�wmk�"���	�Q�,�gN��L�Owh�g��h��?\#��d�=#�G�L=\'b�d�=�����L�/��|i���xŠ*2CN���R���=��:5�k��V�.���������s�ӳ�N�ĽJ�,̸W��:��1:=�UG�'%z�&MKDcf6���hOJ}|սJ�K��ו[�Za_���Uim�o��J|g�)^Dd@4��섃1�u���d�M����m�F�p�3jEdԂ�Q��g��H�5��*�(�.�v&Z$�B�&jL�X�֠��5v;��������f��O���|���vs��ݍp廉�8�F8��z���mv=���Ʈi�1�j ��V�5V_�~/�-�m��J���v%�]��_���Uc_wb���K���4��!����/n��;��6�O5��]���rQc��e6�?�V���>^eQ>n�>Z�>�e��r>����4�������{w�Cy�3{�����l`\��Qc�5��vJcoi�M����O9��;���5v���Vv�C���v�a�C�E��Ca����8�P;��W7��5��+;�ǁ����_c��c����ll�����=Z\#���vk�7N�Kc/�hS^�a/��;�=�N��}��Z�v�a���v��Jc��:(�yl��ve[�����̶j�9,�ƶ��͛"����6b��؆g)4�,|��C��E���a�����8y�ƞ���x�[��@k��jH�:����4�䱕P��0����kl�ƞ���%e�Ɩ8ؓ{Bc�;��3�b�-��>�@Y����Al����y���Y���*�������r��U�+��2N���/4V����L�l+-顔f���Xc�İ�+�a��ٌC�@c���X�� %WcӉ]��r46McS56e�E�bc�ɧ�Cxy(�M�0xtv ����ש�2.�ei,Sc{pK��� ���1��2Fc����lTJ�2j K�TR�Ȥ@e��F�mDK�[�!��ѐ8�Op(Ýlx�g����K�����lJ�?�����7̪��X\]��aV�2�ʆ�Ѹ�<y�� �fC4v���P��<6辎ʠ�l���	Ph��h�/���o4�G_��``���C�}YtG�ZT �4�S"�>m�>�O�ė��;��6,���A��+L魱^�+���b��롱��ga���$�͟�j,��_	�XWW����ÂG� ���.��v�X'X�S�Qc4�����>��k�Gi���ؕ�}X�����6̉�N�9 �#�ٱ������mV�ߟ�뺳�����t��Aw~f��헭&f�5P�h�I�3�cF;3hLiUcJ c�����G�b�#vF�hޒU���=?����?]�Cf��.�4���<%-D�����?�����?��� �;I��:5����?����l�+Z� s�3װ��jv�|�;�'���f�K? ]�g���y��~�Qv�e�FPBv�=��(�,#%<�P���b��?XGv�2�9gO������W� ��+����N���p��5�yd��]�R�����[���T�G�F�P�K�Au?$ d:٪�W6q}�y^��B��uj�!Rp���}R���O���d��	]"�ʳ��F"ln��*�� ��J֨t�<M��\>i�<��"W@s:������Qp�	�/e(iJd.�n��5:V��O�6����ёr2��Ge~��Nx\\��c�2�J��GY�6����+�%Е��&�Y��@��E�J������Jw� ��j�Be�u�Ǔ<�"��F�	ܷ�N������՟��n������Z(��J֩῵ۭ��H�%��v1�V��N��d��Ȓ*�F���)�RM���=��Q�7�N�Jwi�Y���=)8�_�J���s�$�l��z�����PMU�m��}h�Կ�s �^��Kj7�_�Qu^������د���FOփ�d���k�t�b$�����1�t��s������It��Yꪳ^��ڐ���ͯ.�7qסy�3V"=�H�$S"�ϝ��]�v�y����;0�
��߸u!| �%څ��N����Pz���ާ�K���� ���Hd�L���da	�Ɠ�CC��#W�*��U��K�_ɩ�knU��ב��ɹ1Ⱥ1pC��nm�:�]I������ (�د�ҥx���a�7�(%G)Qj�!�e�2GY��at�4���)��a�a�a�a�a��d,+�5��L%S�Ti�y�e�F�I��6y��M�f�f�f�f�fy��L_�^f/�/+/�/^6�lz����(9J�JG�Q��rT=j8j<j:j>jI�!f<K���Te�:�0�8���!B���~�ƴk�����	�vg���.u8T�Я��>v��KV�\�j�ʕ����w��Ǎ�Ձ����J[�����i�,���@]���k�ks�2�](�50�N$r2lg&�ql�,mT��F�1Tb��F<� s�o,l*�X_�������t@é]rujݨ��wAw�¾�Ƀq=I�0EU;td�;����`w��1`�L6J�n��9�}��u�bo�Zǎ9��=�8�k������~0������ �����CCTC���o��l�VK{����y��=t�|�[9�P�ļA�w����:o������/��kӎU��M����d�m���y�i��F5x�kg獡��m_�ٮa���A,$8�����s�`�Y��z����hD�Ȱb��A`o x�M��L3㺭�߾��ጂ7��ܷoӖ-+�>�t�¹��\��r���g��[x����۰���;�T>ڣ�A��?<�C�3~~�e�����L��a�/�0�a�B�2��I�QV���l���sCx��/�s��g�m(��!&ڕ�u�m�_���gZO�Q�o�z��Ƨ�.cj�C�J�rݭ���`�.䁸�Х�F�c�}u�F?i#Y�ٰ+���A�B��A��'=���G_�Ip�vup�����⸾ޕn4��=!�2�k_�s�i����C/<���K{��]��^��r�)澽�k���A�8H���PCp�����v�od;���6�7���p��ڙ�	���R�m���aN��6�����A7ԅ�H�ƴ�!jۀv:��a��{3zW������:���kY�~��˖)��u�>�������o�k7i5}�Σ�����q�w�ݳW쟕�'��*��A	����dENP�Q��jOCH����Aԍz�F�ebt����d���@26�WΏ��X��?�z:I�7�D��qa�V����1��F'�o�����z���o
j�)��w����ݸ6����C7>*�Ķ��0�gtCK� S*|jݳK��{V;����g߻����4��%ͽm̢��-|t�"鍍+Vl�X�|SV�����޾���v=�����ޮ}�N���cs�-Z���BȔ,d�F�i����~c�[i]m��n�!dsX���S�5�7�zX�{���V��y��?���펃����-.e-^��|�n�7�������׵�hKY/m�q9�M��y�P���&m�V�=�U�D��rw��t�󓶓��vU�]d���������rw�=m�8zAc���t4b"aqm��U�k�]�mf2�B]T32�.h��,���n6��%�'yԻ�b������}/����ʳ�{]㜊,Q��=�oT"=����b��oԷm����T�۰�e|��ܕ���N�B��۹]��4y.���*תR-1*T�dLS���>
�xN���$�n)a���r��#q�qmՍ�ed��J�Mc��d�v���o�����ఇwu�qX�'u���}�m7��G��D�K{o��t$�����(m����<ݤȄ	��y�Sϸv*?�n�g���>�Y_+��?_O��&xy��j̒V7VHGf������+����٠m"���xh˿�R�~f��.�/��+��q�����9ő�
z�Ao.�Yɒ�#B�7a3��I�h�� 1bdd�E1q7V̪*G�U�+��]Q𶓨y����I�=���)y8��b4���@��h
�=Y���i �V��L6�̐´��.� ��,AB��?��ܬ}w�Q�u��ҽ����?���.�{�
���K�L��3������QZIz���y<��v!�q����e�7���gו��]j�qn���r�Y�&�d���^pW�1z�u�ҍ��X����#:�Ktp�+�ktH-���R��ֲ�]m�����m�Po���#�?�l����d���p�IG�կ�o�C_}���/�͙��']�nʱ�
e�|�p�������ڸxg��׷:�e����w�ȈY���:d��-Ȃ,*:�c���j�M5m7���\�t���j��.�-&FO�D0s��b���3K����q��e�-Y�b��%���x����+��YW'E}x���.^��dd#}���7�	���U���'��@��:ZW�������a����c�������x�v����0�JlC���9�դ6�Z��	��[�R�=�ۃ�vO�?�wo:� ��x=>���~q�P��G��,�u�($�c�-�Ƹ�v�>���D�F8���\/��-��#����[��>��TW�9�W�9��E�_�d�ʕK�,c�I��U�*s���E 8A�|x���\����?Iq���W��P�Ə�ޡ����]���nj����N��������.qg�߸
_�FW�~�z5t7���:�'�XIщ����u����O/[��.M���rj��W������8��7���w+��Dw���٩�x@�5�^���R1)���%����f�Q.��C�!g
�w�"!)��Oy��{�c�bma�v��~��j��g�i�b�I�ۣ���H��ٳ#�w�u�nbΕmڙj����3�� �=���ށ�����u$6�I���&��7���U�����&@jN�|�۾_6��O�^�l�SuW���3sz��g�El*9��7'�7D�I����w����/ZC�N"#��5.�2��R5�����6�_'����@���߶�8�X�C�U�(?�jI�{Ql�!�ވ���:��AB����_,^YWwߋ��yI:�8J:�q�+�i|Jh�1-���}X/뙐�G�u0 ֓���qU: �TU�T2�l��`�e��4�!/N���8�C)�ђ�RZ�}A����iQkְi�.W-�1��X%<���0����T�$K����pF?X��-s?�������M����A�3��n����s�ٿ�z���������]���'�%O{Q���	؇#���'�8Yk�������?�9��Λ��Z}��Ra�ڵ5�֮]u�7��r�&���?�����j�k_j_h�>47�H��m���uy<�׹)�m�'��.�E#DT���馐�$�'F��ݳ_}����^>]��^{J��O�j|[5�ɜ���}�0����'t_�3��'�����&Fl����?1:��N��L�;����0;�S��E\��&H�ю8G����$����·���m�^~��y)��ϣO$���F���L��Of/���
~���8?�d��2�$��}PpPB��@�%(XnKV�cr�ʶ�krM���]̖�N2��jK1�!I=��p��o��k����^�"�����B�N�`q1W}�Q�����4�6s���_�|U���f�8�5o�wƤm�\8=i�<xd䃙�G��:n]��Ph���s'.�O��[����
Y���������m�џ z�x�l��$8��ike�o9)>փ����b9��]�2���/���ì�v|Mc����v�Q�����͝�)���f3=n��l6��k��c<{�������u��?���W�{��_�/��Ʒ�4���/��}��32���pGȏ�3ׄ�TR��I�8�'DM@�y\Q�u�)$� �b����U���k���4m��ˌ��Ha��sʾ&�b�Q�D��jG�b�������x�RG\����d����L�Imo00i48VmO�	fEbF�����b6�Y`1��3zR�x�▜�9��S|r��I��`�E��:��ΦN掖`k8A�,�+=՞�Pc�u�4@�6�5�&SLɖQ���l��Dk�T�
�"e�)�2K���1�7UX���;H�,D�����Roe�4Tbi�h�))��G��l��P���7/4Bo���(���Zh����~�v{����gK	�G���k���-�]S��%Х��7Ri�T�=����H�Y{�),�1���d��a1C����-�2�����I)F5Ɋ��p�sϸ������/�F�LT5�"�,:נ(x1�5���̓��f#d4I�&���"���֝��W��:���I���/7��׵a�H)P{�>��Z����:Im\�_{�w�d����8�;�����N��a���������m���Tc8�o����bp�)��6���(v�����U|�i�brR�p\G�>�.Fgk�p[�� G�#�9���0y*�6��8�K��&rDnH���K�<B{���'ha�Q�VlZږ)'崆��X�U���DB��$<I��C��s��>���|2o� ��P��r��@Z\� S;�i;`Vjd�$yN~�|�nU;�d?����j��֑����D>d�z�5��z�'w"��?����5y���ҿ/��la]����c�uuZX��o#�t^�2��ﷳ�|�N��_[�j78��|�Ȑ��[���d@�2YHC��~I�[��&��f�8͹��y �^d�a�':/��W3�|8	o��>P%��q��5�E?�"���֑�b;d�\(�����_P(yJM��iP%���A6�j�q�9��>6~l��RM ���̫�oZ��}������oރ{p��=���܃{p��=���܃{p��=�?���M�����@iGmMa*��UJ�x���IY�_;hn�}�
��JO]%6��S���v��n!]�󞺟iy�S��~hg��&�1�{ꔸ,���D���:�i�}�
	����U�ْ�I�e��n!��_y�~m­&O�F
-�^V>��hFa��GnOWLtt_�������ʪ����WJin�+��ؕ�GU�2�+�+f��E��g振v���ȯt�T今J]��Ӌ�r]ye%9E��1�9���1e�e	ee��ϯ�,*+u�D����n��]PV����|aUUylTT�gUGV�UW���U�ȏ,ͯ��]�HQTQi^������Ԣ�����d1�s�%j��գ2?�5=��lv�H���=�ln��s\:�&�����������j�"�說���/ɩx�UVК�ٜ�_QRT)�х��XkFENiU~^����c��"\Ue��ҹ�r�ʦWA��X%L�U��C��斕�c8PU�ź�]=B�JBz�X�+���,�(�A���%��U9U����b��(&�2�
�fC�!='��eyչ��L^+�^]�/xh1!V�-����.�*,��3%E����
]� []��\�WI��Zط�0�g��fTY��2v��"����Ҝ9�-犮�N,4�����	���X0_L�+sU�E�*����ϭ�-����\�ܲҼ".Ge�ٜ����e���	�����
f��[�Uʛ=@�sU�@�����8yN9�J���������[�_���"u�Z������K��
����W��Pќ�<!��:��r*�WuqN�X(/��hF�`cF����J>�{hN.�T�^~*[��{\����b��x�yyi�K�纊Z�:D�����!��J%W&��w�����uf�U�U�B��b_���
�[7D���D'���ĩV�\�YeEM��ϩ®q唗c��L/�������0�9U�JP�/m�,���y�j�H����q%D���,[YV�w�07T���G�����Grf@0��Ҳ������RZ`1���352ɕ<6-˕969kB|F�+%ӕ�1v|JbR�+$>�!�	)Y#ǎ�raDF|Z�D��dW|�D�蔴�WRvzFRf�kl�+eLzjJ�R҆��KLI�J����Y�Ԕ1)Y �5VL��JI����$e�����Ԕ���䔬4N3D�]��Y)�ǥ�g���e���L�D�MKIK��*Ic� �>1#e�ȬL�Bc�++#>1iL|����X���C"�%h����ə#�SS]	)Y�YI�c�X��ic�p�KK��J��JH�(�	�I:oexj|ʘWb���I�͋�aq���'�HJKʈO�pe�'O��1%#ix�	�C����c�2����.��LK@�x�7\p&�O���N�،�&V&�d&E��3R29�c�.�'fp�A��xi~��x۝ށQ|�G�Ĥ�T��l�1ޕ4'7�����gs��Q�R=~F�Ճ \xD)6��&��g�,q���ys�#9�~y��w�4��oެ|D�JJ�?�x0�]T)v:���2ϹW�S��0�i�eN1�U6��rCy��"L�]QT�`�ʩFkE�<�Q\�9�ZK�Wi�E~e9N��Y��s#1���g���Rda%х�r�b�1��5Cσ���"]f2�t9�K*H�A
Iq�$���3�D��6#\$c��XWat>�!%$�)��#��5\$��V�x��3sf�a��$�6Ɠj����P�!F�P��]�R
\�1�A��\�_�usD_k:��
�0�JQP��#���WbV��.���-�{g{綤] Zu��<�s	��_��Ӥy��0>���_	��V�"A#s��l��J���ϝ��r�,G[��6_�O�}����k�;m��*���vˇ�ʰZOa��5z�~�n+�z�A͗�;}�,�<�
|��~��	��<Zt��a���G�V?�)^�d�^����:�Bї�k�X�T�c��S z�V�-��^��LpX*�{v�����*����W��z4�Y%�h�#rė_p)�P�R�uދ[�4�V�����刽�_�Q)�p�|���+K�*���O������h�y8�U�����u�[ʁ˰J�೙�<!A������5~x��^�gՂ�����
E���h�D��J�_��+un��#|���%^[7��J̎�9"��Q�%(��A�]��jK����^��ܖ7ytU+�k�h��G��Z��
D�-�H��b��|��䚘����>�׏�=Q�k�\�v����i�؝Y�Y9�X&"C�|cQ���t����c�{���1�w�KȜ�������5]z$��{����}�x����c�
~D�#[h���r��m�D�"�����^�zz��)�i���}��{~�Ut}U�J���(Op��U꣍��}�)\ٴ�7����}׻Fk�T��L�1.����ݍ���z��r7#<v/�~$�Wx"P�௤]oKe�gz�M�S$���[X`��*O��˹�$w�|�����6}虜:g��}_��k�g?x-1�Ew��ɪ<g]�O�Y�f��_���wL���.���/<��E��n1��V{�H_}��h���鞭��{f7�:��DqSR�ђb���G�gx,����B����/"�K5ݳG�<�bA��F�$��X��7��X�e�	�'3D���.�s��7����]�E��q��X2N��id s���i��;��i���&�?m�W�TǢ�i�Ak*�I�q|��qx���g��zi��%���y�9�B{�-�J+z9�����_�*hM�'�zZ��Nㅎ8eNs88Jo�u���)�/dֹM2$�_�%Ip�[B�h��"��b�s�Y��R�gd���˓(��UG�V���+�z3�H�.u>���7��)�O���Yh���}/]���4��8!_���X�B���Z��Lm��c��B_�n��D�R��H�]%�Rki��y�w�B�$��T1:zL�����S���=��i�~��D��v��eĪI���k)��C8��R�����>:k�~�ǺÛl=VxٝZ� �b�/l�٤�d��x8��a^;�����&�Z�׻���~N��iy�ni�D�O�3����t�ؕ�s-W�w�s�ǿ�'�o�؜����9��fz!Ɩ��ܪ�g��j����pw;���d=�o�~�ه����o��'�t=�l�J��)3�-z��t�6X"F���*ź�d՞�i��e���j�w�揝P�o����W�-�U�̄�W���絺W��U�������+��ˉ~�*��d��n��Ϛu�5�V�����ǩŒ�y(����<�?W�k�� ~܏�����CH�H�wN��VaCy��ށ0�)B�e�fԶH[PN��ۥ_��Cz���]��Fz���^�'���A��Ko����ꧤS��-?J�<_~�0y��.�g峨�'�����a��P�����eB�{���Z�.e����L��[DMLN�"�99�It�܊b2tFE�#$�8��E&�T��+M�ſ��k�А��̌�0�Q�
���w��1%s���-p��cƦ��:�L����ɱhi���_����+y��[Q5=O|S��5�"$T�AHi����lG�H��Ƣ�p-��l�o5�52<�9�������S�E7������Zt>��N��M�B�頥xv�J	�U�J南�ly����L�'
��	��ќw̑r!���o�������"�	�������Q�3��t�I�|���I�Aڑ��b�]N��琞����D�����}�G�q/Øt��M-/b�Q�jl��垆k�Б��h�c�I%B�����Qk	��|�ᘡ�4h���s�5����-�I�d��R;��"��"�~R�'%K�R��-M��R�4K�/=���ZZ��Y+�vK��:�tR:-��>�.J_J�����6#LeV�d�,�uc�X4���6���,6�Mc��U�9�1�$[�ֲl+��^d{�~v�co�3�}�1��]b߰k�&k�%�(�� �����9F$��Qr�<^�,O��R�J��/�k�g�M���y��W> ��˧�w�s��s�k�^�.ߒ5EV̊]i�tVB�J��O�U�d%U�P��)J�2S)Wf)�Ǖe�je��E�Uv*��}J�rD9��V�**�/���U�r[%��ZU�����^j�:@�&�#�45K��NS�b�B��>�>��Pתԭ�v�Eu��_=�S�TϨ������o�k�M�� ��!����2�"1�A���D�(C�a�a2l�-,�����4�����h����IU�l/��g�o5���
��=_�>��s���T�Z�Ixa�"�KCԥY�r�b���Ԗ	j�D�w"p-����C=@���C��y���w��Jq�~�ź>|J�/s�>�y�+k�_E/��-�H1&�G���׃ࡿ���,�����i�\*j|8Y�	����'p�hyP�l�+p�h�&��r�������*�%E�	�%K`}d?�G���9��3]��!z�sL?w^&��>]�*��d��n�G�l��D�H����G�l���A�/��NhI_(���������ݱ4Lp�����A���]��։�]�Tn�I�b���kL�c88?�8нH�����z]+�,p�V#8�8�kR*F��b���'�6�7���G��,w0i\ۄ�b�X���T����E�|N�&�u߾+���ީi|�������p�fzÊTh�N֠j���u<G�ki�V���g��1�&��>�����zaS���5��&��{���^ժ��6Ѯ�>�:�h�]��L�b>W��q���8�]�u�F����+~�ow?,,X�vM�Ԟ�A�9���	��m����』7�������F�'ep��e���GJ���yo�`��=�H�i�?���p+H��J>KC!��L�9�����Oę$i�!8[=�G����	H��F���2����X�H����7���o��̶&X��9�d�.2Ϻ�g~!~��W~=�z�+~��"�7��I��e���\f��-��пU�C��Z�3�l�ST���[��L�˿�2Y�l-͹�	����=.?!?)/A���p8ѿ�.e�P���(��\Ǔ�ݝx�-�2n��d��g�ӗ�Mz��O?���K�z�ޤ�$%� u�\R�!�H���R�4JJ��K���R�T*UI�E�R�FzF�$=���.�NH��㸇�#��.H�K_K��u閤1�����c�Y��"Y?��X2Ke,�Mayl&+g��|�8[�V��l�e;�n��ձ#�$;�β�E�%�̮��LdU��N9P��ɽ�hy�<DN�G�ir�<I�&��r�<^���B^+o������=�~��|L~S>#�/,*_�����7�ER��M	P:*.%\�Pb�A�P%Q��+���t�P)U��y�"e�R�<�lR�Wv(�����r\9����S.(�+_+��u喢��jV�j;����P#�~j��&��j���NQ�ԙj�:K��>�.SW���-j��Sݭ�S��#�I��zV�P��~�^V��7��bP�T�$�x�g�1����n=#�q{��t�x�k��s��x�ސy�e���H����)|Lᙃ�g�M2�I��5�/*�O�(�~2Ɠ�*�^=�#�҃����,��s�U���k
r$�V=)��#o�<�^㔥*���ny���T:,#���
�;��ci*�nc\�"��d�'��%�	��8V���	�8�WJ�!��$%���_��/sʢ%K�T�K��[��ӵ
�e�|�kU��'�hw	[�KM��E��|uzP�݂�lQ�'�N����}�+�"|�����'�ۥ2y��!�s�|Th���*����O%�j��k��ɷ�Vwx��%/�bZ'�vQ?��K��e����
��yޒm�'E����ܣ�"��#�����q�J�.��OW9�B�}�.񺕝��Ux��s
h��en�������k�2?\J��ӄ�q��qo�U�çq�e�M-�xL���Z����y���3�Le~�Y�݂.��kR
���o<��x�^�$/~��w�_�g���-{Cx5�A�+<���Ϊ����� =�6�<����i��2��t�;����x���F���N�(��~��ǋ�5�Ur�>@�T��/r
���*�.�j���g��T����n�����n�K]�t��D�z�&��o�!�4D5�lG�?���?�bV�e�~N�v���<��~�aܚs���b��K\{�)��-(##B����o�6�6��E4��x����~?뉖>��xS�[Z.�[OO�©	�z,���c?��q/�O�<S���0�I�a&#�a��_�Pܨ_ �D>�C�3y"�)�L�u�5��X����L��_w�3��|�3��|���7u3b��z+�H�R��M�%EK�!R�4RJ���I�4�@*�*�9�cғ�
i��A�*m�^��H���қ��}�c�S��tM�)50��?m,�ud.�"XĆ�D6����l2��
Y)�b��"��հg�&�<��v��� ;̎�S�v�]`���Y=��n1M�e�l��ɝ���)��c�89YN�3�ly��'ϔ��Y����2y��^�"��;���>�N>"��O�g����e��|C��EU��S	T��nJ/%Z�Q��J���LR�)J�R��QS�TV(k��Ve��GٯT�)o*g�����O�K�7�5�ҠJ�Q��jGե��j�:H�&���tu�:Y����j�:O]�.Uk�g�M���u��W=�V����w�s��s�k�^���R5�l0�v�ΆCC���!�gH6�2ن)�<�LC�a������[����݆}�:��I�i�YÇ���/�W7��Ĩ�F�1�d�f�e�601&Gӌ�r�O6�{��Q�'�cE���Sʾ�)Z<s�zg1�R�ګ��b�;0[w�}�7}Z���g�Rа?��u_�&z�1!��I�}�t��sL}V�Ƿ୲�7}��D?�u�����u���~>4��i����GW���ȧЪ/�ա�����?Z�Z���<�~N}K�w�`]��/���[���!(�z�g���u�s<������y�9�x|�����/��n�sg��X��~��_��D��c��Հ;�����Q4D��>�~@�-�Q�ξvl���K`��l����:�gj������;|=D���s���x�gh0�~0�s��IG�8y��#+�&K��H
�E��r�'�$y���S�_���Ϥ�\$_a��`�u�-y��$�$�m�@67U�Vj�m�ڎ�'/ӎ4�����P�
�}ɫt }��E��^'������s�9J-/X^���%�K�Y�Z�R��{�~�X�Y�S��S�g��_�Tz��7m�T�!�c����鵟�;�tC���Pe�gXdXj�1<c�dxްð˰�p�p�p�p������s�׆z�u�-�f��f������b�a�4�3����Tc�1�8Řg�i,7�2�7>n\F�q5�z�c�q�q�q���x�x�x�x�����K�e�U��m1�&��i
4���z��MLCL	���4S!�I(�P
P�Q*P�3=iZ�i-���(�Q^Dك���	�b:�o3}��)
|����&���%��ن`�hv����p��p��p��p��532\s�y�y�y:_��3��T� ��,E�Aye��(;Pv��E9�r�|�|
�wPΡ\@��ks��:��P4B,2��bn�׳`�YBPz�D��ĴĢġ$��Z2,ٖ)�<�g����t��O,��,��*���v��e'�n�}(u(������b"��C���/-�-W-7P�M�}V\���X�(�� >������'��u�5x$J�v��iVX�*�L�v�α>f}Һºֺ��պ�
�Ya;�~�A�cb�g����[?�~j�d��k(������`;?�_�_G?�n'���?XΏ�M�_��(?�L���&��z~�~��_������r~5���������]~��l�w�8
�����n~�����5J�,�wK̇�l��Q���`=lg��l�����v�X[�-ٖj˰eۦ��l3m�Y����m�l�m�m[l����ݶ}�:��I�i�Yۇ���/m�mWm7l�����o�w���w����?����H�4�,�I������+���?����
������o����~�������?��������_������M��d7�m� {G��n����ه�����������B{���>ϾȾ�^cƾ���}�}�}�����������9����������[v�!;������#������u�9���G�c�#�1�Q���xܱ̱ڱޱ�Q�������sq�t�v�u|����q�q�q�q�I����t:�A�n�^�h� �g�s�3͙���,p;+�s��9������*�*~��xi�p?n D���"d�W @iS�c���@�UT�@S��Ҵ�)�Ц��1� ��"H�vF1"FDZ)m<��n�웗�?�̹��ٻ��{νw�����mF��˨7�M�A�q�x�8a�6�5��K��q���8��i�If�9�|�L5'��f�9��2s�<��\j����Js��ɬ2�͝f��`6��f��f5��'�3�Y��nv�W���M+h�[}-a%[����hk�5њjͲ�1fe#-@�GB��{-�^��B��{-U-�_��B��{-�^��B��{-�^�����k��Z�!�:Ϻ�t	��B/��Rm�b��6�~�@{�=�c�ٓ���l�{��k؋�R��^k���go���5�.���k7�����-��}�~�>g_�/�W�k���8�[X"I��HA*�b�Hb��9"O���L��b��$�D��)�D�h͢U����8)Έ��h⪸.n&��&������ÝY?�Ν��[;��4��z����z�#\�*�F��W'�kc����"'&��{�[���ύ�-~�+<|W���R�Ꚍ�N���S�:Dǎ|/�z/=����u��U��{�F��~,���1K�q+�shQl����=n˷T--�[��|{��L��Ůbz?�k��黺��ܗ��^_��Z�����3>8�Juj�:��:�����>����)����w������s6-v;����{{�^���:�}��rT�E+��,~u~<��/ʌ��2���_[��P�O}���&q@�����Y,�Y�ov�.�k�w���$������n��3]�A��}�w��j3~�ؽn�+�ζU�|�� ��m,�:=�S]�(�Ө�k=ur	S�;/�:�:��M���=}����_F��o5B�$g�]L����y&���Yή$�n�����[	�ҷ�A�{=4��)�j�{��i���B#\L��#�f�^���Z��k��Z����u§[��?��	'��om�����!tm#�F�*_��B8ű�鄓�~���~�U�n�����NO�/ߧ����h��BWdIw�N��i��L�a,�dL@6�l�3	�$�O8�p9�r��o�v�%G�m��O!<�p!�B��rT�I8�� �b�6M��\MdJ!qJB2����x�'�Dyz���"�������!��w���΃��s��#�#��R��$g�Ds=���yzyY��,�'���лvv�q��b�����1v��b�eW�Z����Ɨ����$�v��'�����-���h&���$>QKצ�"-C�͗��������<�d`�<�Ϋ��|K(1�ȷ���F�gBCyC�P�9���{�U�*�Jxkx+��o���5��*�����y����̛i���-8��I?�[%�mx�a��b��eP�Vm���Rv�`��EYc)�C~���HDzI�^D������I��3�d �C��c��I�c�pM�'!M�H�=�$#zre\�I���a����zჴI�8� Ɉ�z��$c��#�� �O�N�2^��u��vo��gP:��Yޭ-�c�O�����/�V��|����2F���i�ԁ�D�J��mbU����5�F��ZY��qv��ag�y��:Џ���<��y_.x2̇��|�ȧ�Y|��x>/�󕼂�?�ȷ������W��w<%�B�����	��r���2~�3�����#�������e\2ʵ�GH&�Ǵ������$߬�K�)ã��Dڀ$��d4`5�>��~�ƚ�KGW��
.�r�Rtŝ��U_��}^�qD��L���Y��YDy�e���V�漓�r�,�(����4:35�|O�zu�	��,�Ϙ6?�e�|,��i󰤼�\�ͥ��\�]Ly������Bs)/4�d�~�N�������OW���Z�ҋ���d%��%l��HY!ˊ�EV�d���ťx�\�|QI���˚��zw��ݻ-���ւ��������~L���1l��f���K]I��<湿˘N�c}�9ʑ��(�Z�{����q����~�dNE/0��\f�Z,��!T{����汇;�@f/��8�=�4�������/���v��`[����6e��1A1���I9���]~��m����& �IV��0��4�3a<��W૰����@��rx�O�:�߇�O��?��a7��`?����[���w�?�?�>A|������p?��/������J4�r\�����F&������a�	�c�5�:|�a��5�m�.<?��Vx~
������u��}�o�?���a��~� �"���5��1 ��G�,��FP���X`}����@=^d��/�\W�Y0�!r!��ʡ*a=<�`3l�j��Z��z�C�I�X�����k�e��^��&$�@������l����che�!�si��s4��ZC�z3���S��ɝgޤ3-t� ��#%�<��hd�:{T�3٨��9Ԃ���흖���H�� �X1ۨ�y��NL���<��舾�qD��Ɩ��
endstream
endobj
20 0 obj
<<
/Filter /FlateDecode
/Length 421
>>
stream
H�\�ێ�0�_e.�+b|�J�6�H��AM� ��1�!y��?�EE���y��f�����Q��o�a�s�n�=5AN��EQ��]3.*�k=H1���m�C<���J�cڼ��!O�m
���ڐ�x��_�㤏�a��!�����6����������������<1�"~>� e�j�ѷ�6�MHu��n����~z*	��o�8�ӹ�]���y)7y�|B}D�P/yQ��o(���*Q{gj eP ʢ �C(�P�� 
@�� �5�µ^\cW(�j �]�[_�(9ژ������e8Cav�ƝZ�\����!�0�s �R�b�R�b�R�b���+��p�XLxJ���K)���X�z|Z�z KZ`��,>=�Œ�M�t�ܮ�T��BsOi�<z�����bx�Ρf*� `L�P
endstream
endobj
25 0 obj
<<
/Filter /FlateDecode
/Length 14941
/Length1 35396
/Type /Stream
>>
stream
x��}xTյ��g�s&�B!�W	B��~���$$�2�LH �ę�����R�R�)E�Q���R����-Zk�U���"ZK-Er���뜙L��������b���~����k���r�q�X ���M+�x����5�����O�N�Hc�6�M�K��~��?��!T/�^67��i1�0v���aY��ݽ�1���Uջg�H�c�h��U+�\�
�؀�hsku����F�_�X_�Z�42�Վ½��nu��}�[�X�v�xݞ(�����S�����ϸ��~@M}Ӫ_<���Sp��:_�������|��ֻW5�ժ�~�����<~f�mq�/�\Ϯ��	����m,�����;G�R�9��ȍ���<�o�o��7�r6t�P������֪��sԛ}@����9��D)���,K'֥ q,[Rc\����<�4ƴ�ڏp�l]��X����h����~�҂o�|BrYIu����+����Q�?\�����i��Y�}��?dc�ݬK���h����e|(�]ǮgO� [˪�&v���g>�,�
�g:��e[ٝl/;̚q���q=�汕lۅtz-d��x�2�PF��aװ�]�vX%zo�})�[��#�c;Y	ڏeA� �������c�'YJ������rCy/���-P��}|<�e���6`�b��m`$CV�C
���M�b�/�r��$CrYHa�DH6�^Nr��t't��$Վ��"ӝ��`i�C
�cј�Mhw p#R��,2���ȶ#T�S$�sp�@����L17���]*�O���Co�t�I/��Bf)5��=�07ɹ��au������d%��d�R�l}X���7��Ǻ?<�B�-�&�~�b �� ]��9�� K�K}Iy/����,1h������$�MTڃ�6���>>{�|���(2Mf_�F��\���Г�h��/Iò��vIjt����Y��y�7�jdf��x�g@o���g�iX9���`U��7�xv�F6� �2��u~����KX������'AI����~���0�J*�\VN+v�e������0z���� Y�38�	)zc���氙lz���l� p;��̣���g�A���]�>�}��P��P�x:���.�o�=Ю��O7_�}�@>�s�����a����m��=�b�B��1�3v/�z�_��}�/��;����_�y|"_�˔a�A�woB�%�^��Q_��O��S�<z�3�k���Ř�'��!ׯ�����������xC��g�������f\�fK~�0�^�ȝ�����~�u�ݝ��JXS�0Q��hƲB�n�f+q/��e�� ���Z��+1����,�eS�J�l��jY�9��`n�1O��`�ð�*X�jE����U���m�t������[��g�d	(i���}?���B�Nȭ4c���n+F����t^VH@�P�X�*=�ȮB�X�#� �G>b?q��Z[t���{z��}l���-���;�&x��(9 :�C4���0�CN^;a��K��T�&y�J{�n�~<�^�Kw"Or�V����oi�c�F�;!����6(E�9FopJ�F�Hy�b��N��t��;]%Vn#�䗁n�>(��(e!�B�l��j�3�占8��bem��l�TD%%�-��r�/� ֕��0ڭ�jߋ1���=܁�ܟD�� ��~�M3h�A�J6�e��R&dt�/���^��}�a�H��-D�eG!��O�/&'������f?�о��$�a���pv�F��%]�8~��A[S0��Ak _,?¶`�^`�ZAc��т�n�����3��Om�>����l4�i�����_5�e1R_P6K�/l��qѼ�GO�ο���<�h�=�����eG;連.𩽨ă}�X	���W���G�lܕ���ao՘�X�M�a��Y��3x`0��K��{�.�y4՛�n���ߩ�7`  >7�w�A�)u��lDYw��EMwV�'����:�ff�n �
i "��*�e���<�����Zo������3�C
�%K�R(��"#��X�Q�B���֬E�R�X
��4�"b*Jr�J/(ES離�KET�1G�i_��#}�L2.���d��Pv���5�R�쑱���"�[�S�Ɋ�4�t��u[�f�:st�<����=�p��/�|��֚�1�UYnG�����Z.ll�hU�A� XU,�����7��G^h��f�s͹�uep�N\����zk���_h�p���r� �L}�2��/�k�wɫ��7<�(Ү���2~�,�i�6��6�|���Qt�)}�\��t��~f��]~��uRO�7��L7'�YX- y�bQ��7��V���W�sb����X�o��\���jh8��Ea��A����l;�g��v�;��cq��^�w��qfd��{p�K�݀�D�ƾ�K��)�A�(� u�����qM��i��q�!�_���a�H��(Cd�E�@>�%�4+m)�x5ۈ�D�{������щ�8#?�ώq������pO\�w��;�O�sYAD]n8��`<�%vK��D�E��5=V��sVk�jP#��mGW���~�ڈ���9H��}eе=U�Z�~�QVB�������T��<�Y7�]����`	#5�8��a��6N���g�s��a���`~��9��-d�Y��=;��T>�^�����E��)B�{S_�?���"h�v��	�c��tB%�kE&%�u�	-��Nuv��?t�	�/ӟ�Oe��Zp�#v˅��v y�8��9m+i�1�%>���i*g����S�ů�!�V[9��� 9����`���ǚ���]Fm�W~�`�?Q��}��c��=�8��?��tր�紒�_���yU�$�/�z�ͥ�C*�����|����и��_J��$���2�VCt�tyPj-<�N�w�5ħ~	� W�u,_��LB�%��|,]�%���h��7�Sl�0@�Ys4���	��M��Έn��{'�G��}n�.#O]��[���v#�m���F��.A<�f/��&�d)j{�U����۱��v��nXg��
��O�F�Ql2����������g4⬵�����p�Y�V�uL�-Y��N\G�T�G$������Xp�	J�p�c�Sf��<+?|e"���6�3A"��8%�ǉ�+����b0�C���D�� >G�:�]��
���4%[�c=��-8�e�������F�?����z¿A�A�m�� P�c@a8x�ޮ/� ܍ �����$}�+�Κ�S��'RP����P:D��_�s���7a_AKAvt�؁Fз$ռ�O�o ^f���z���Di(v�2�1�e��� DJ���y��*9����d�f��`�Ѱ�4�~Q�.�Y3Og��h$��.<��=����D~�(�#�v��w������<H���
9ؿ+��<
���*B^g�.��|�W�OgO @�?�7��ǐ�\���?��*a��2?�^���z��iu�W��/w�)w�L8�J?|2|�|(� �t�]�ς��+��)�����v���D$��q�~��#��|���{[��� tّy��j�w���I�9�۾���������X��{��VNt�kX/���ː����g����6�TN�/	�\�~<�����6�o��ދ�j}G�>�Ň8y(�'v]��C�v>q�Y��]8^ݰ��$��� 99�?g�Ӑ�|����iN�r�Z�*|���C����Kx�Rk1��i�W���US��[5�/�n}.z���1�7�� )��([I�<�NÑ����>���HӐ��IF�v*$�XI��g�R$��d�\�vZ w��Vr���t����E|s�Y_����Sc���ߡM�}��>�Y"e����u6����}~��5U(�e��*����s*\/,�74�í+��:�JvZ�:�T�����Ej�A5���o�<14cVI���3�y6��%y(+�@Vޡ��yT'=���_������]qw��pW�w�PvDY��t�O=%�|J<q^��8��t��S����P�x�E<�%�-��]����]����!S��y'm�y��Nb����������ڃŃ��=?K��,{�՟��ݦ�i���M<�s���)8|=;���I��s��I����,m�r��,�����΋�bk��Tђ$�o�-���)6�b�7N۴V�{O�vo��gc�vO��'�N���w��Oiw�b���O���;nO��X,��VoO���Y��������E�l����>K������#n�*nlk=�2q=(^�%֠��,�:I�B�*�Xi��h
t�����L�o��2E#j�
_�h�Jk0E}�b��)Q�N��M����lu�r�7˞���TQ�>5���Q�����7NxLQe�JS�׊%���#]��-2��	ba�X0��� QT$����6���\S��9��8Q��s��1�$N��(J�D�)�f{��1�#
M1�3�j3[DAW1㼘~^L[+��j�kE^W15I�Ċ��Ĕx1yR�6��&:�I�b�SL�]��"Əsj㻋���qN1.[;&I;V�sc���QI��Yb��mT�� �F$iY1�#���aIى��<1,Id�(3Y͈׆vC�(���jƐ�ZF��8�0���,����n������u����YbPg1p�H���������I��H靠�d�~�QZ�)r�(ѷW�ַ�H�%�}ФO�� z����E��h�g�x�gW���GTg�G��!y��&%��D"�%��ncE�Xѕ'k]ϋ.Y">.K�?/�P�%:�Vh�׊X��V�N �)Y�Κ�,��Eʣ��YDY: ��)a��kњ#�#<���E�g�=T�E��&���,X��p�m��!��?l��ܧ����v��gx[Į@�@�HQl�j��87,�[-b+��iԍD]�:I�V�(���&�!N�z�-^�P��&�ee�րS��h� ��=8==���,OE��<����#~Sp}����R����0Z�f����uP��{��`o�3�[�V��-�vW��я�	�����γy��������`G�je�򼺄�z�8�,R�W�������'`�[�6�9�څ�,ƪ��{�����`���c��bojo)�q~��b���)����c�ˇ9n�Πw��p����j��Fۍ���zf�Q��QZ���aǎ��⎟>~zx��~����ը�B@���'��{�K�.����b��z�h85��b��F���K�qv�KY�9hH�q�k}K"�y��׃��^Ȏ������jrL*��)����㻏���11�`�6lҩ�c(��Ł���(<;�#N��#N����)�n��|qvi��ѽ��J�2Y�*��;�u�Î�c~��ULlw�t1L��9g��J�����&qG�����'⾨��w�Į��я�_��QOF�\��:S^��uPúq�t�׋���/�������G��?�4!�uʦ�C���垯�)�4�����;?�n��a/���n�F��=���ѣr�9��PMU��<��ݳ��lub��t��:�&�N���5�`c��=��,9��Ξ>{:��Wg�����.��e%v����S�n	�#�ƌUSg�4[��x,��Q�m�6ͽ/w��!|O������ٱ��{h�+/a�q8s����z�j	�gMlBM�?�N�$��,QɊOt���)�����>%���2�,��R���.#�9�3zTx�� �a?�>s�w�Y���Qw��^['�U��qz�����I�7����ȑ]H��E�k-VS�O����n��f�6u��a�E�{�HM��%2#36�W���ܝ�p�V�鸏�ĝ!�g;_5^��j��^�-�od���/�K�	ңC-�>�����O��?x��h��G�c��)�F�*�����[�]����ٕ��<�*^۴����2+��O'�
���a�N(�k�t��&������͝��'=�K4��艮�t0}��iܱS��))v<TK:�����R��Ǔy�����'��/��E��<����-.��+��[��ɓG���Jn��~������Ϳ~ޫ7�|��"��9�㸅���m*�}=�f����nFL�&�YW6�T���q���t�؅IǤ1����
3��c���7%��]Px�y�����%֟8�����Z1�4�^'���EcQ|�h���V�!�]86~��c<�'$N�rJI㷘�S�J+?5��~��)����W�6�xǒ����8Yw�?��^Ӎ�t���?):�K�H4ғȚ-k�;3�����qı�)L��]��v٪U��y������g>3?�<�=!���w���Ϳ ��Ǟ�ԛ�vӳbDtK5�w�c:E'2g7HvZ.#}�X���,����j�6��yUo�~��Ӓ���C]9)0J��ș�V��zA]r`Im�ޤ���w��~�=����:�&GE+���ɩ�1j�3��ʻݝ�:�&��ߨ5�w��%G;��r�)�c�:RF��"�p���H�/-9%��[�9�%�����!.���������tg���)=6�밄a�2�{��ION���o��n�y�u�U�y��ش1à�ѣ�@��9WTz�v���������ݿ�f�Y��ٻ������:9�F�?�$K$��|�/~ѿ?gc'L?nRJ��]v���0#��+����":����f�԰I&�u�M�{β��$̐ms�l�����G�M����'���y����gf�x�]E=��`���^]�tV����@S5�k��T�r��`�9θ�%�1�{���SY����e'��*t��%
m���0M����b��@���ͱ�zqu�������������Xx-bYhM�ݰ��By���ƌ����M�E�=E��+!.M�ʻZ��ϊ�/�SƘ��f�K�5��`5�fٽ��T����o���I�s>�<��|��q>%y�-p�;���d��?ǟS�E������E�p���W�
\�+p���W�
\�+p���W�
����+p.��'�ǆ���,�?n9�Ý�W�3[y����Ո���d�u֕���Q,�}��;Y���w��>{��ǲQL��F��h�r;ϙ˙n��e�.W#�Kr��y��9Ct�X��{v��&8�󝺦��|,�q>6�׸�_����5�*ݕ5|�HW�jWnmS���u�g�
�2]9uu�R�*�*���^OfL�w�{^����ݰ�p��^Wm����������ջkBm���l_�ϕ�������WV�ȱVY/���j�O���5������	ÆyP��93�k�Wy�}����oӰ���k��6x��2k��Vy�i�[�$�
���z]��:���L�w� 3&��3w�,�a����'&�װ��ȵ`���w{��n�r���#������6@�E��ߋ����M^O�����C{�&��ݰ�Ո�@_e�mX�Q���l�T�'�]U�oDs٠���,M���JR�A��r��Z7ƃ���M�&�Oumt<HR��2_u�J�<%�8�{�>Os���xj!Xmes��xh�!�TU�쑜��m��57���Z{ ��o�d�h/��p�{Ij��@MF�r�a>�+��<�u-X���0�dd���l��@+k|�w��P��o��^����W��r���I�X:��IJ��|�Z)G`BLL9�ܕ�^���"b l�&LC�*����fV�+P�P�^[k`F�n'��v�w����K��jZ��vc�L������Ւ~��S[]+�]��CD�In�N�/�|5׹�4���]�@l,�[�X������@$ {��	tɲ8��0w]�D�~!^�(�ņ�ծ�v���^��7j+3�L97�%��y-V����+%�S�ء
W�\�)�6̎��V��ڌy�B��Ն�jªq���ܕu^Ya��&����q@���^/���=�f�H����~%Œ�r3�[�ʦ���v�I��j��Z�^
����C��V�������Z25#�5����UV<�|~Ni����URZ<� /?ϕ�S��������s�]hQ�ST��U<͕S��5��(/Õ_QR�_V�*.u�.),�GYA��¹yE�]��WT\�*,�]P�����&U�_&���/�:�9���2\�
ʋ$�i ��*�)-/�:�0��U2����,4�@���hZ)Fɟ�!@hjqɂ҂�3�3Щ���Ҝ���9��2$����EM2�%h�����e3r
]��e��9�e[���Eų������r�!JNna��D�Z�S0;Õ�3;gz~Y� ��-N�:d���E��9������2=��O-���=4QH�N-.*˟3h2#��� 9�7�8#� ��S^\Zfe~AY~�+���L�0�����D)�\�SN^�ͯ�#Yv�u���m���S�e����º�WUy��mۋ�r��J-��AVk9���,\����g�,�y,׶�䖜a�_�>`�؍,��Y�HW����dem�V:��z����u�­�/�u���~A�6�F-����6�����(�׮��b��Uu�@�ґ�7Ј��v��nu&���~F��6 
��E'�U5M��&�R"����2]1l*�!�^����-e5�]l�b�f�ထ�U����M ���^2���ր�����E�Xi�V�z�{�2��!��f��B[7�,��.�%}�4 7��{�pW�;��GYבNQ�f�U��ه�����GT���H6��P�P����ǩ�zK�&[R�&�:��L�c�_���h�������O�f����z%�Z�4���}W��4QVH�{�3/�1vHO���x~d]���ZΡ���s%�������Lz9ץF�4�F.���-��P��9�����E�Z[�.�wӬ֓V���;�6^�d%D����ٮE��꼶\Ki��Gѩ�Zox4k�-�� �|�a�o�ׇ5�T���%��d��5��D\�_n��"i���(���u�lZ�VJ����̹i-�k���B�-�e�U��z��D5!�T�1[v<(�c��SH���,;�#��D�4�0J3��ƍ�$h"[�/m����<B�����Y3Q�t��l��<D���z*��(D���*-n�I��#��4���n[����92�r#/�"��z�h��Zm?���:�9��ưE7u��6�V�>����PM����1���#����JX/$j
����:�K�f����ǵ6�hu�۽��|��� ��i�bO�@�o��@�����xI��E2�홪�퐭Yڰ<��2���e�}=]���ٖmV���$��v��\_���a��i���Zy4�{�����S7���m�#�.��Q,}5�����$��r�"���^�(w�@x��u��X���~�*S���07�ѥ8�<'��먗K�a�{����W���K�շ�*	�-3�n:�"^��y���J��C�S.�/�����C��)�f����L%�{_���z��
��^Bc2&k��ٺ`�bn��p����x����!O�k���K���bIw).k��(2R_)��WR���?�fv��%	��Њ�D]8��=�Sl$�^�Ԟ1k_���������f�*�5�d��aM�*�q�Y��8Ÿ+g�O�R�|ё�^t^� ��G��C5�>�V�|�%�bz�˦Q
,i/@���{y7�@K��g4F>�PI�,%ڳQZ�k��N������{���d4j�W�^�vd?ɋ�i9��Fm�U��l6�JA�]��DO�A����0��lNsHG���9ҝ,��k	ڕ�>sHf��"�a�-Y�k&,���Z��e��r�B�Tn�� 	�<y�_�:�J-Ί�Y��6*��.->\�:���H��:]$9J�inr@?D7d;Ӊ���%�rH�4B.�I-J}�[�F��Tҗ�7�y��C)��$!j�g�R�a:ɗO�*��e�c>��K,{, Y�ں�hZvo�Da�v���rf�`�|ۦrHw�V��M
krl<5Bgm�_d����\��]�����U�uYX�h�ζ9�aa�y�k�gq������P���;,Z����`�S��aYX�N��]��ת�c�k���߹#�Ƕ�42��`m�62���tj[ߡ][�埭=����]j�
�����-�E���F�ѯ��t+��k���#��T۶�[��zjy�и�d�v������Mт-p	m^n��xBl���e%���D��l���k:���NU�6!Y�M�~��Ff��jI�2�̴��Y�|֦�뻰���f}���1�:X��Ǟq�{59f��v4|�7қ�/��2�E1%�ߘ˘�>7�ufB��qe��#�)ې�_�1�;��WoP�`Bݠ���k�kȿ������ȟp�d����S�22n<ba���W��2�]cr�v�}���i��,��wW��U��ul�R�w9+�s�\lQ���JSI� �o+�����a��4�DF�G�8��Q,��l����E�����B�"����٨�YeSI�X��$�F8�~y�r�c(�C���)L���d�r�%g4K`�� L�(6	�.H'�3�k���a�%�7[�����]$�ji�'��}o�����+�Z�}��	���,�G>�%Gkɩ!�$�ߖ:RoVo�U�7���[Ȇ�]�_��)[�s���(_��G0��=JQ�d���7�����<.Y<
//�F湲=�;\rC��&�u]�$!�%�Z+.C��p奠�eY"#	oT�CGI�m]!���W��Z_��~�����芡tQ��de�2X��Q&)���H)W*K�j�N�+���[����J��]٥�U(��'�g�_+/)o(�(TN)�*_(_)�"�D�H=�K���%Ɖ)"O�%b�X$*E�hMb�X'n��U���>qPO����q\�+>���KqN���ƨqj��[MQ���(u���NS�R�B�F����FuV��X������ԝ�u���zD=�S_�*[}O=�~��QϪ�5����EKҒ��`m�6F���j3�"�\[�-Ѫ�:ͯ��n�n���6k-�vm��W;�ҞԞ�~��������Q;�}�}�}�]�=J�����KO�3�,}�>E��g�%�<}�^���z��F_�߮oԷ�[��n}�~P?�?�?��������?�?�O�_��tӡ:bq�DGoG�c�#�1�1����(t�:*�8<�e�F�
���g���R��B���E&�]�� ��
�I��@��z�z�P���pF�_���3I֚��>�|]pk+��_�qE����E>��l�B�{�|X�W�PKp�!� �j`��W����>�����PI���ӭ���T���cp~*\�Q���Δt�r�;h�"���U�5�pq�\CW��nne��V�cJZ�u�٭����;�Z�h�d�����(�:x?���v�˒�󩤜��r�YT�Xb~<�Y�����R�<���q�[啄����.k[�KYպ�t�Z�|���fm�=������A�N"��k�A%��X�q)��#>��g�����?�ޡ�<�	a~�-��,�C4��.�k	�fN���� ���<�xs"Z.6���|�4��0~ ��k.�sM���%��	�?���3��/x��F��e1��a��yp����r� x7�����s�+�Si���՗į�~~�@+���(,&�#*y�������oA���7�6�M�n*�ʟ�%wt�9Ĺ��Q>"�<��?Z�cw�A�t��rFz����H��G�Z�[�,��/���!򿠖�}�k�,�s:07�I��7X,k�V���b*�.5F+�kJ����W�?�6�I'HW?��Z�����c���H�`�Kk���גg�$K��$Z/τ�?+�P�by�����Aʮ�4��x�(4b�Q��r]Mq��Y
bLi�7Ҙ�H72X��dLb+���=W2N���3����d߷#�W.�l�et�cn��M��%U��J�G��P��o�tI[d�}|-�o7������!V���7�YoK��2i
R�ޡ+{g��\uI�%��c������f�*w�;�����Og������(J��$(=���d(Y�8e����TJ�y�"�R�Q�&e��N�]٨lQ�*;���>�rXyZyNyAyE9���|�|��V�T�)�PE�����H�D�%&�l1M�RQ!��L4��q�� ���mb��#��G�qT/�����=qR|"Έ���T]5�.j���P���1�$5W�����Bu�Z�֩~u,�V�.u�ڢnWw�{��!�I����K��;��S���W�MѢ�X-A멹�4-C���iS�<m�V���i�Z�֠5ik�u���Fm��Uۡ���i�����s��+�q�]��#���vN3uU����D�����3�Q�=[���z�~��ї��
��f}�~�~��Mߩ�����G���1�E�5�m�=����~F?��w0��0]I�d� �`�p��$G�c���Q�X�X�v�9��U��:�rlv�8���{h���hw˼�ų�kCye�(C�+�܉z�r��R�
�G]�oȾV^�a���
��?R�s�,�S ?�;�o��Q�g�ԟ�c鈔�a�+�_��T
ɉ_î��,�H�U��2",k��w𷅌�V9J�*[�W�J��T�G(�b*є2M�nP���V�j=�'i�GO��+q����E�ܗ�'��Ϗ���&\��&<�p.�%��Qe4U�Jyq8A���Z��ƚ�Ӯ��I�\�-����j8�(��
�p�㣴s�㴗�W9dT�������Q�b��CF�i�.�!b��}�:UFz�ޢƅ�o%��Gպp��D��2���Z.?���r!��|L�^&W����/��I֪a�c����s5D��Y�	*9+�#JJ��a�ۖ�U��)�r��oS��iQO/����B�a�&m&V����N��Z�Ԓ&�Z�-w菑�I
=ɮK��L!��4��Y[��U�n�Ց���9a��}��x検G~R�3?��V�*�w��p�*��+�~m��y�zQx������m�u�%�K��J鲤}b]�Q��tpF�.��oP���"�_GdB��Iq�F]�C8S�}
�e
�����O��y��It�'��P>�����!�{:�cvB����%'��>�>��ه��T.W��bc%Fr˟Ԧ�t��[1G��p��G��d�1W�L3��<�y�-�r������P�HM�s��1(y�Z�$<��1������Y��,ii��,���"�BI����B����2�xx���G�|����r��/&
��!R�ʛDM��W�L���G}8�K�Dm��}���s��uy�����ˉO�pQ>����W_B��#��j EP�)���"�f��VW�l���8�F��>�8����(C}Mz�D72��<���D���A<���x6��y)���p_��
~��o�����6��������?ʏ��k�m�����t�5f!�~+�#<���;o�hSsQ�ŵ�1ߡ�%�K$��Qy,"�4"�f���s�5�\}�<Q�)]d�H�P�P���|.��~~�?��H��r��@������3�	�+�8��N{��D貝�9��C#'ص /�:�o��]�L�dNlEl1�:�x���#��rF��Fs�wbc䋛�8��s��=��u�:��?����/�K6��o,����Y��32��3�q�'�a��l�X-�e����>��]l�c�c#�ulrlb�[��刉[X�s�s/�9�9b��_8��΃�GX�y��8kv��|��t���[-��NOW=W�º�odlR%R���h����uH�#mD���"���H���#=���H��'m�?�qrV��N� +N��(S�;�;O���w;d��v@�}��0dyr��w��#v;Ϲ�����!���L�%�M���?J������p��u��oj�]ʿ)9���+�>��LO�z���g���|�o�Lz�/��in�4g��_&˧T���%�^[�|옿=k���{֘E��ѳ�
z�XI��"��=m��|z�����v����W��Ss�]�$��xzN!0=���'�����@V��
zYIO +�	dE�I'sd�p���NFW�^6�SW��M��mp��چ�&6nVR竪c�/��zjY�_��a���~fi�C�%u���w肰v��V�����z�ٷ��ZW��~�'|�z�Kc�S��η��|B��I�4��B~�׈8u��m�y�4c�Qh���<c�q�QiT5�2��h0��
c�q�q�q�q�q���h1�;�]�c���8�<������S�W�3F���F#�Ht�FO#�`6R��۫�֙��؃����g�g�\���F�QnT��%��h4��U��:�Vc����l�gl5�;���^c�q�y�y�������0��8#�`Fo�e�!�VX��Q0S�Q���.�YQk��C~�:�k�G"��ɒԟ�o?m>���2c�q�q�Qe����Ҹ޸ɸŸø��d|���q���ƃ�@�a��ο:?v���w���p���Π���k�C�)>8K�K�d��)�L��s
��NB�@�����Q�g<�m<<%\s�jQͣT�F�'Y.}*��+v~\H[������K��U���ö����]���ϥ�Y�����L�
endstream
endobj
28 0 obj
<<
/Filter /FlateDecode
/Length 281
>>
stream
H�\��j� �_e����n�B`IYȡ4�$:�
��1��}�	[���ϙ��3��}i���>�z���:�0�4�3�J���)���n[<έT���\���p�f�`�N�Sz��w��VkpF��uǐ起o��������W~;�_��f����F�b{���Bu
���V��?h$ɆQ�z�󬎆_�ɋd�G��('z"�D"
��g"JV�%�
]r��{Y�WR=N�J��)YY�F�ǖ�����saT�{Ҍ�t���Zc�*�_ Dg�
endstream
endobj
29 0 obj
<<
/Filter /FlateDecode
/Length 2878
>>
stream
H��W�n���W輀i�M�I�0 )�!� �-�=d�A|���!,�8"[]lvw����!M{f��X���7)f� �O�i��S�������������\|�WyTVH�+�O��}�������D��~~���������/&�^�}�R{)�$����QJ�⫍?2?k�,�o��w���i��g�/�����9���Ɩ篯������X\%�y0�ك�����9��g��"L���0u�IC���_c���I-"��/p�����5�����|�L=�o�������#@v�\#�Ą���V������H��i�B$�&��/x^�d�]���2=�jpy@�q,u�`��ķFx���l�� ol�̷��3�u�F*`(���g����9,:nO��MB%).e���f3T�kw���L>י��ӼA'�9!Y�̰֒m�t���,�Z:�%񄖼H<��k���'���Z���
���[׿t5	�82D(��tu����l�+��<WJ�oYئ��U��HJF��d��"��*WW���ΖFۡ�7�Iv���\W���P�1����N�;�yݿ���.�r���,�7:Oq6k��~��nS�� gS�O4�yH<��;Μ��q(��q �8~cFQ��q�@~:<��l~��h���ya ��t-��#k��K�u;c� ]`}rY��x#F�6u�u�����[6�?��$.(�;�D��9�X.��ib�6�ύU�-��M����gK�c{����!|�����}�L�T�[/7:z�wQ�
|��N�j#������Dw�ܞxdЊ@l5-��AF�����VП�<87��:�����.F���j�mSѪuNH�*!T��c���t�(m!�)S������-��!6���KZ�i|�ۓ˽u	8�aJoXzM�2�/�C��(Q�:���4W�b�W��/1����y�,w��}��u�U��{ޯ� �����~|g�S�Q�6)ߓ����Nq�z���Yc%T]c4�8�;�pg/_��oV�-F�t-��0
8=0�xb�5@b�IS�)HE���?��0i���X
4̼5��5c�|8;�;��♙I l#�M/�N"�f��e����p�E~:n��|���}��0�iO^���<�Ϙ�?��y��`�j�s�6s����8ӳw�a�1LsUg>3u�g>/[`Ǚ�zQA����>t{!�=m[���Ũ^�ł?�ŻQ��b+��j�0������z����ƣ��M�n�����	�>i�
��:h����*��Ij���<U�P�#C�<E�:]�y�|�SP��i�!p����(���bz����Sz�l:'�g������D�N��X%D!���� ��y�GE�Y�C!ƿ��2����@2 (V�2uuMd͠�)B�����t�E4�LM�څ�3O��߲�>9��[��Nz�� ����=}����n��j�2��˟h��G*[o�c��`�:��GG�Q�M�f��1��Z�L��]������v���ٹ�a����\)C�a�6��y��k\�,�\��)E �<�J�Fp�����l�3�V˄��K%��Q��{��D�hz�_]ߤ�U�_h7�`ի8�XK�D�9� }���Fё�&%&�o&=��xeAJ{����i$��{��$�D(� �N2��@�&O$�I
����(�����Cռ��y9P)�u1�&K����8��B���5�;K�[���ms�V57-;[�qFLL^��9d�F͏�;	�T��?F�kP�~׎���bY�_���"��J��E(��J�����=�]������~AC��q҂�$�-7	�m2�eA8�Z�����S,�ib}�diӂp_�mq
܍� ��m���LFLL�
�2l��M�Ma�\l�G�c5z޴ ����샸�2�`��Qh:E�'��@"?m�D��#4��O����?�����z����i�o,a��[Ǳ���L�ӷ�#t�)�M}�Xc�Z�<eND�`��������sŠO�� ��1o��ӆ�'&W�����+FMb{��&��M&�V�+F�+*hc�8O��$��dis��*�,ڲ	p7��6�}+wf2�`b�.��!�6j�\1�I 젚���9c�Fϛ+�ezF�A=�2�|Wu�h�@p�[1YY1����?�����X���}`f��c�����w���{sŸ�VL�+�T*��c�J�c����w�!�`�`�]pg;�rjp��η��8�x���1֘'�q��\�JTFhJ:�����Y�i�k�l�9�s���j��P;hqڦ>�'�ǹ�����c����-XW]P�é��㨏Dؚ�!'��"t�q��6���h<��#��y)���6�[oX���v�p�W���E��S��[n�۷��iI67夸��3�`b���q�!�6j&��rA� 젚��1r�X���,��T>�g��s�+�UF,�8
M�h�o%B#�]k�����%L��~c	sL�:�U��d
옾u�3O�n���7if4�S��C�
��[�`�Jv�`a�^)pp\�0஼3�LL��aUC����v4'���8�j4nhf��������ƿ�ر��d�S;E{^�%�a�O�3��[+��	�y�kvL��6�VS`�t>�D��c�F���!�3�{�L�b0BS�Q�o%�^�rN	�b���9c���Hk���6'L���p��V���b�4����kj�׭D�7f����H~�w8�/����
�\P� R�� O�K�69z����7l����טԃ�7]�y�3	��3d�厨U���b-L^�S�A���H���  =�-�
endstream
endobj
3 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 4 0 R
/C2_0 13 0 R
/C2_1 21 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents 29 0 R
/Parent 2 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [3 0 R]
/Count 1
>>
endobj
33 0 obj
<<
/Count 1
/First 30 0 R
/Last 30 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/Outlines 33 0 R
>>
endobj
32 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227162914Z)
>>
endobj
8 0 obj
<<
/Type /ObjStm
/N 19
/First 141
/Filter /FlateDecode
/Length 2598
>>
stream
x��Zko���_1c�� V?�:M-�."�c�Y$��}Ϲw�\����)`��rw�s�cfT�5ͤf�	��d���D$)�4�j^�֌˦D[��H=҆48�)�9㽩!!H�7>"-����!-L���Ԅ�P���}��Ͼ�n6��������������f���h6������|6�<y��y�7g���/�������R���;�n���z��l�1�b|��sq�b�������f�K�z��͟].>ܚa}�9=]�ǜ�xt�_1�Y�~~����D?^��V�+����Q�au��9m�o~X|\��Oyr�������~��|�\�h����r��3�a}�qq�/�jO�E�^n��wO�>\.1���f��Bz���3;s��ެQ翺Q�P�Y9]�.��XW8[�oQ�˫�M�1<}��c�]��٧�7�fvh�_��[sn�y�Xy,��J�:�ZAI��#k�	1��&U�&໤�I_�>0?���z����`2���I�dRF>�o�wf����%��!�Ao z��&�A�X�ɮ���ӊ��. �cI賦	���#��f1~�7y����1�(�z�9�G+�+�m�8�|�\�r�Ơn���kB������-��\� ��%潟�<�|���r3��?}�\���O�k̏��}C����� �>`�Z�l��q�������*� 8��L���%Nrt��N_`�J��{Y'�e��Ӆ�ʲ�j�]�^Hr�)a�z��2	#d@����8�$B�a�-AF IH�!� I�%1��瘗C��>����c����
�wْp��	�-���
'.��)I���͙��+SA�B�g�m��lż�����X,z�tȆ"�R����W,8�H�0��5�|$M�<�W���V�R;� LO��<�D��XI�,�i�)��E�M�%yi͒j;4_�}�$*ꃯdݜ����O�0/���#&�~��Ry�%��s�I���k�������@Rc<bUi�Y$x��{���%��l�.}�A~':zG�ML6;Vb1h"L`l����)L-�A�%v�%�i�{�SВX��hf���`*���	+&U�/�`<�rF�="9���]�;��G�C���uδ���,��Ј��3�lC��T����4��J�&2�����!�j�
�t7������z�Ǹ�n��S��*�~0	����Vj3c�K�/��b�M}�~�����`<2�66A�1��e�A3�.�b讚X�t]'H�q�6��"le�BCl�\���[}�3tx��a߆�#�}D�Ycl��!h���j��v��{N�3=uq�%�����Q�[��9`"w���_8���a��n�� ��#�0�iGQ�3�C�%�����L��_���k�qt��Cv�o{�;���铇�?����~��4�o2�@ܡ���RYk�;�d�X�
��|��S{3�K���vJM��KHm�{+�}$ٴ��lZ��:�,�j�2�2�Ü݇C�Y�=6a�\�}�y�[ێ�z �y��;���H��pۉ�Bo�+�Ɲ�R�.('��0VI�g�iNhKQ"�WX�%�����
a��i*�c@D)$Vc�&�8�"�u����\�m9�R	��,SH2�OҮ�E.�mJY[%�Ot�)H��@v1���j���w҆G!m �>���)�U�8�����g�θ�$��C���z��l<�;=/2��v_�C
�R�N��UJ��R�θF���;���8�OT� �G!t0))��SSR��#(*c��w�1�P�ƿ  (E���J �P���ն�J����2l�8��@&t�y9`���C2:��}�O� &v�kߪX쇜���ws��Z�,W�~�E��]�$9ۺ�5V��2 d���2��$��/���Q�9~�cVq *� ���~�~�{}�gz�/��X��O��G<�G?���1Д��3�t}�7�|9��U�t���!��ᾈ��0�G�Ǣ�#F{5@_�?8��O��N����lÝ���u~�]�>�ػ��[]��P�=��N��^��*�e���T�W��r���w������7�\�P1_\���<��bt��W߿~~z�Lo�/�6�yk�^t}�n��7���F��������Z��j��K*H��M:3���/1�O�(OxjK��z1�0;G@.o0i�IJ�_�#R�#R�#R�C��[V%�G$yD
|D�|DJ|D��J��S�����#fm*�� �H�V��К�q��\(�H	m����]�R�AS��I�x���:���U�[E�x�/R�яJ��G��G��G$1�T����Ȫ��Z%n����i̽���g�.�Χ��_��ݒ��d�ސ��_��_���7��/��Z\�|�rwx�����yk��s���Ź˻�oވKG7�Ñ���G
4���P]=��ճ�{�Ǐ/�\����*�#�=���Yw=N̞����'�?J8�G�����1�|�$�� �Ͽ�|���C���7������3a�e��y�y���?���j����ONa�ͣ�����/��o���r]�
endstream
endobj
34 0 obj
<<
/Size 35
/Root 1 0 R
/Info 32 0 R
/ID [<51888BEFF55B2B4F9AE414499E1C2ADE> <C8662BE9F20DA503331D56BC1BCFC9DD>]
/Type /XRef
/W [1 2 2]
/Filter /FlateDecode
/Index [0 35]
/Length 122
>>
stream
x�%α�`�;@Q!qw!4�0��ha�oM#�0�c໼�K�.yy ֕�	0�����"���n| QY�`�w{�[�cy�!ۯǣ�E!Jv���fG?�jqbX�Zo���]
endstream
endobj
startxref
47549
%%EOF
