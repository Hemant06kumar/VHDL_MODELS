%PDF-1.7
%����
10 0 obj
<<
/Filter /FlateDecode
/Length 22
>>
stream
H�:��"������� ` 
endstream
endobj
11 0 obj
<<
/Filter /FlateDecode
/Length 2248
/Subtype /CIDFontType0C
>>
stream
H�|TyTS�~1&7V��&��V*��}���Ȣ�� @X�0	�
�B$+�"�P��[��R:�Stt�LG�::����}���/L��9=������~����w�l���`|�us̎���R���m��c%�y�b�7���S�F5�A͜J	|x�<����q���g��K�@���8-�'c�16���3|�6��ɒ�T�L)U���Eriz�R�x���^\<�K&1l�O��%�����d�D��DqE
�$G!�����\R.VJR�6dg�&K+Dr�B"��N�܎H�I���\$���RZ/����rq�$G,����Ѵ���H*ѵD;dR/�Sғ
�X�BW!'WI!�dJ�T�X�).�(W"Z!J������`�F�a<����~�-a+�O�MX$��`q�l'��I�����z��b���c>�fʜ)}�y̛S���� k5�4۟��~
�g�W��2h�ʤ�=�nԊ	�Cv��Y�s����^��28ɐ�Q^�ͤ�+�{n0��	�<T�.�g�B6���:�P�5��p�P��>NPM >o{aT)G	.W�.T�u	���u�P� x�0x�
��ݏ��^��7L�� 8�[��pHX"��0Z �]`�Mo%����;��}��g�*6�T���͸�2!�
�e)���6EW��q�[і%<�Y��r��t)ڳ����Kȅ��^��iğP�?0�����C�]������ڥZz�2 }l�B�p��3�C�ʸ���V�B'��hJ��t��&��8-���C*�E᣽g�(l)�O7f�x �5v��ao��!;���c��ϧ��2^IJ��P�`�^�ߝq��PXT�m `�w�M^'��2���z1!,`���:%x�wi��uy5y��N�L�5�X;�e�=$�Rc7,&<s�*��s<���A���W�n����A��������W�Q��Xl)�?�x�����]��L�[�_����*�,��d�(���Q@1J���T�ݯ�ЈJc4��w���Vq��w��9��x�UņJ�)V3��,3��Ypt�^�J�!	��y���`@���/�����d�kQYS9�l�8�X��}��Q�¥X�ۭn��Ւ�����д��o'	�����wF[._7=�� ���:or	,�m���.���\���X���k�|p�#ڄM6eC�����?{�=��Iwr�։��^?�H0�����ܓ�(��?*�<⬪�m��$�����\dO������P`B�"��?�I�Kb��IE`�]W�8�u�����#�/~ܞ|"SSM[���F��1��~I�K�3�P��)�;���^��/��J3k,�	�H+�r$A�Q�q��A��h6�{�J����1���n|T벶�	�{Y� '�Z��k5s�^r�W�H?�Ώ�8�ù��]:�8�!�JTc0���a�q�=O���;�4]r8���ڛ0�R���5�&N��bo&��rEܤdA�>��Mb�������������ĄJa�V[$�������p��%>%��ڂ�o���܍��T7����:��J�*�rr
�	�y�yNe�X���_��d��n�v�IM�d�Y�ݪ\�ftNl,`<u3ay�W���!��@��>���5#:�a3�����#�&]�oo3��a�7L����s���q��^���6WD�]^I����km��
�i\e����ӿ��ď�SU�++���]��]�{ß�+.|�Tr�-O�1:�����
�^��a���� $��W�Qs���ڢ� P
��h��]�CN�Ϊ�{�;a���u��?^�=R/ć����Z�Du]s3A[&M<�;G�EKT��]�^��;Y�be��/�l�Jk�jm���b�Y�����$�+3����5=)#���Ս�j$=���kk*�=���MT�YŒT�mW	���v�&���?^f���dJ%G���8�	!pӘq�tJ�K,O���f�����6�<�j�7v
�m�mMm������/��p����í�/K@���F<�΀�R8I��9o������y3����6�s�{���,��� o����Jr����ykyjwlwnP�y�������\r���Z��n^pcoh�cY��M�q�O�W�������������	�p��`�q 
�&�	[|��I����%���������F�_	��
��w�c ��D
endstream
endobj
12 0 obj
<<
/Filter /FlateDecode
/Length 287
>>
stream
H�\��j�0��z�=&� ۱CƐ&-����li�
jY���o_y7�P��3hG�T�kk�?���j��8{����X�f��
7��Z'd47�p�m?����)�6G=v���k��^as95[����h$PU���A��{kI�]��n²������!d�)_F�'�*����(�x*(_�Z�O������w�i<��I�%�3ә(͈�)S��3=1�2�rֲS�ę9g�Y+X�?2=�r���'-r��Rl�}���X=u��c,�_Ѝ�k�į  .��
endstream
endobj
17 0 obj
<<
/Filter /FlateDecode
/Length 23026
/Length1 50268
/Type /Stream
>>
stream
x��	\G�0\Ww� � x! �D　�P���
��Q�x$Q�F��7�u�5�!j�(5&�D��11���,1�1�5��=U��c�{�����O�z����箧z�A!��!K||����B��
������������p�wpJrZ�����#����1㖯Y���@p�FV�/߇��Gff��\��1���t_��rˍ*ńP����ܒɅc�SW�X`��ə��-��{�����=�⃐�����lņ`<����PC`<Ά�y���̉p�m�)�Y�z"�p�3��xlS���Ka��(�0��_.�!���J���m��XX^R�S��1�o9���VȊ����.[5�����߀�χǻ޳_^ހ�#�~p�=�?0O)Tۃ�.����)��q�"���F�A�
�^�$��!m�[?�J?F��&8�N��a�@!�пt�Sr㲑Yl6�S�ě�B��D��ڮ��/�<�**a8V?�P?b�;�8�e�8�@�h��6�e�Z�h��o�(C�;�-
��+`�I��/CgP!���H譀�
���������o��\<�Zַ�	4�	Q����U���Z���K��	�u�Կ�>	|���lzC��x `tEӀ~��Њ���S�=�^�9�oռ��4xN��^�{Y�k�O�M���/���L�`/ �z��� ˢƺz�2�c�z�!5�E��P4�kYm6[=�� ���r$�qS���:���� ^�5�!����q]!$�T�A7���>��`��fО�� �=�z�/���������-���Q=Q;-�Q$,�;��^P)#�����ZP3Mm��	uDC�&�\m����g�g~=�����m�
�sy�F��F-!г&�F	qlE� !C>� ���ҵvH׊}�2�'$j_�.�9h���Z�.'���w�
�\��h
�8|O�G^�ɗ`V����B�@��1�s�n�3���W��E{a�,��L� l�[�*t
0g@o5Ĕ<(���h��v� %Oꫡp|��n^��F�&�Ά 7�� �W�I>\�2]�u{���?� ��|�7D���h	�}
:]���P���<�#@f����
e<�θ3���g@9 �?{/���x����8�c��	��!^�[�O�? �������7�D�p(�����b���.����$�5�w�1o%� �f7�2��)sf��@+�#�!F��������<��o�?�������@�o����l����%��pow?xl���a#E,��x���
��
��3Ў����=�U���7�X}u(Z�h+���?��F&�Ѡ�x1k���F�%(��x'_mz�?B�B�����1�g[����@�\4�+�Hk;��6��B�w(z8�<��v�_ �t��/8���=%� w)p_
��wRđD�9��`s��c�k(u`�_'u_��,;�s ���qIh�� �|i�ؓ��=p��,0���1�|���%�c�?����<��J�h���^%���G�	j���,�h�>ST;�6:�-"�
ASS�9=Ѣ�����y@ko��6桮p�bÓз��	p	�
u"�Lų ��Z�_����g}�g�/���a�����6��C;���`��a�&�<ۂ��� ���nÌ`)oBlȃ@���(�	�6ؽ�C^��!��xF�M�՗� }5N�B���sP:@1�̠)#�H�:�ЃB����}��bJx8��2�q=�b1h�,\����ƽa��a�8����!�< VC��>څ���8*@3 ���2Q����4LD�,(9P��$���x��F�~8������P�V �MGq�[�44'�n�j��%����K���-�������>b�K0�%��x�ZS��
x���j�_ �{��
�X
V2j=����%G�V�C��mq(a��1����Ł�ƃ�t��e0N�}!򎅙P��g8�l���@����,���e@���y� ��g�p&`�B�����`�(p����pt[ �s���w��}�g�jϪ�u�~u̬n�{Fe�� �e�g���Տ��R ����2��b�Q�l����R6����XJ?�	?��c�</h�g��8Op�q��
{u�Mxf�X��<�r�ZF���2j�@-���)��l�E���\�܆+TCÝ�|X/���V(�֨Yj�_o�~�q+�A���m��\u���!�^f;��}I]Q�YQo �8է%�0'W�y]���o�/�H�_@F�[`�!v�����7x�]k7�n[+O� � �p�+!�~�q��C~ћ�+F�~�����Y��@�WN�X�!����p�j\Q���v�{h(d�?���܍m��Vdak�<��^`��a7�����h���m�<����0��J ܿ#NjC�	�%@�1���D�J4�hg��?����;���<�<b��<v4~�+�E�.�0v�0�ý���<�0��W��G�t(C��8;�a�s�q�O�M��@On�Xk�e4��g�hm��^���S+!�>%z�~O��6����E���؊q�+�zi|������ �ЬĈ=X�h^yFy@�D	����h>�gux_�Vzs�v�,�1Q{�ҷ�e>���D��u� �Q���ʨf�P�?�{`�H��z���d��{�,�bo����@I�K˙���||2��=�=�i��td<���>E�R���^I0r�Ff���`W��`�Rn�+��e�A���]�qM��bos��{��6��0�ɶ:я���{�s���[�!��C{�苇�g��V�md�#�/��}����	�@3q����d�r�:�OCn���J|8ħ�sm��������������p�����}x��B|t��(��<���	�z��B�xk�c����S~H�
�.d�-�����K�C��<O��.rF(͞l9����3!���@��@���!>G��Q�¹���0���;g�w8�����yT^\!��j��� ��D3�����z&��0��؍x�9���9(^�]����ٝĪ�p� 8G -}��h���_K�l��Mj֡� �T8]��H8:õ;
å�7NA� �<&��`=����N	� S��]���C	�K*��pV����pjj��!�A�N���@	t����n�A����l���$� 2+����ᬲ��o;��� �`8��u �0�m�� �#a\hE _}`� h{C	�'���kg�m4u��< ������]��?�BT�R�A��Hxn�[8A��>��.z���'�4T.j7��i {�3�DqF�z�d����:�n��s���
�x���rB��'�>+pg�	/Ƌyfd�̋x�v�
�R@�����1�G � ��!��t;�O'�D�������p�Ȱ�p8Ɇ�jI��/���B|�,%�����o&X�7�{.���Zx���ئ8^�I�W�pƝ�+2��~����q�H�k�-<>�Wȣ��jԑP�9���5��|���σ���H�������׵b���A�DPd��Փ�W��<�]g�u��F��۾W��eq���h��;��
�p^����۬(��D�	�5���R!w�/>5��>)y��7�B&�)�f��ܖ��$g�C��`���=P�V���lS�^ ��7�oB��w,���%�IP�'\�"G��I>�X�S��!�bD���3�8b�`���c��q �|��S���gb��x>�#`��(� �'���q�� "�t�m6�׿Q���|��_�1	x�Wڟ3�f8Z�|�����u�9�aP��i!�.��h���v����P�=\���x�j$�4��P{C�W��	z���	���P����K�N�:�t�3��]t�*��g�� ��+����ӻH��[�A���ͤ�<�#숚ݐ�W\���z�~�����v����,��`�! �N �.���l"t� !�>-V�,�K$�4�<�;��D���O�7r���O	���8�ɏ�W�_���^Wd�QȻC-�$8!{�������B[�Z̊e/J��2�Rc��d����R��4ذ�}�K��:,%�R�[���h�&�BgZ4�tC\�x�W�+ÿ��{-Yy����AQ��9Q�� �׾uOJ��l��<İ'R��J@pQ��E�,���U�]��s��] q��fF�3��F��I�2@2G�"ڲ#�6�T�у��U���a�W��*�I�}�ޛC�[)��ҟ���?���Vһ�؏wB�G���N��v���}z;��K��T�}$��I�[O��:����.Xm쟃�7��o�����J��M[�*��-��J�=E�V�W��_�J_ާ_�ҫ���*�L�W>�����S/zy=��'^��T��Jg�/���Q�7���E�~��Q�P����W���ݥ������*=����"XzG�gUzf=�ҷUzJ�'7�H�*=���*}K�� �1Oz�D��yH:��7?)�y��9�>,~���C���J�XOkVGK��� \ܧ\�U�Z6ݗM��J�z�=*ݭZ�U�K��;U��W��H�Õ���]z���N�g[7���m��U�U�/��z��T�M��d���җ��F�Y�/�"/�t�ݸ!Lڨ�a�
֯ZO׿pHZ����^8D_��֭	��=I�Y�Z�>������CtM0]�XMW��<�JgZ	��tmE0]�N��t�J��t�"wi�J�Ӆ*]��g�c�g��|�ΛN�>3G���g��9~t�Jg�ҙ*��ҩ*�(7In��#�eVn���X�-��R�>����I��iQa'�(�v�*}*�NQi~$ͻO'��*�Qi�J�&�IY*����$?��҉*����c�����l:�47c=�g
��IG�t�JG���FD�t���4U�O̡)*M��I*��I�U�x��D�&�HC�ЄAR��#Q�`��M��.����ۇ�q�y�A5�jub1�nR�;��!�R�������:�$Y]��σ��&'i����Vk6{\����i�>։F���_6�۽��w����<��*�5���h#�F{���J#a`�J����mhD�p��-���B[I�<i�5�K��h('w=��%X��.0�K0�L���*�Ҏ*q���1Rp��F�T��&�4��M
�C-ݨ�0�+����Jہl۩�-h��/m�R_����5`hO���I�1���,yu��f�
Ƶ�0�C����{5�
fwj�d��j��ܨ�&;W��j����\@v.F����LN��m�sV�81��ɛ�TQ��e�J��s�>l�$E1��Qd��g/Z������������y݉��k.�=K�\������;p��j�;x>���t��p>X '�2X ��������U���C8�|
��~��Q �
ؖ5�B�g�' ΢Gh�:
�6�0΂5��\W�
��忍��%P֢m�ڜ�@�gh?�]�����ù�$У��+��� K�Kv�$W�n�j��7�p*c�r})]"]�~� �Ih�tI����K�-x�P{�F�T��.���0�N�Ї���N�ѧ�xb���� :N��K�dO�Z	B��\<�Me�Lc�NtpN���>@�����$UJ����\�I�֠lF��� �爊��x:��b���V�O� �i/X�͒Vj��MZI�~!܃�i���@�]�f1��9��n�Ex?Ѝ�9�L�s�'�����,O������<
�1�� 6H�L^{��;2_��X��=�=8�= ���2ڶ���z����R�x@#�t'�
\�!��e-5 Fd���
�t�]dv���}a�t���+��Lw�#���-e0��	wj�4rD����x�z�V���[����EWQ�]a^d�{�~0��.���ӣuP��ӣ�X�`���u�d�k�c��]���&>��U\[x�ގv�
ǫ`g�a΀��.�	oo/O����Փ�qg5`�=���W�T��]ǧ���Oqzת_��8�F>Vg�G�U��G2��9;B/�
߭?�)�����s5^��UZH�l��j�0��
�D� � �M�~"�������	B������9~� |��wW�G�����5Kp��X6Z���q��3U������˯������w ���7a�kw�z�f���p��&��p.���J�!�)��<��@:�������N���Q2N&��d�	h�@&'8oA[���na[�-�e�a����=h�C��=l��Gޣ�1�q�c��|�G�Qz����G����NG�G���}):�M�&��	�	N|�_B��I�$�ٻG�����*���=zDz��IG�D�zx�)���[�rŊ��V�X���?~���;�f���>}��f��zF=����7�#����|�Yu:^���s�o*c�`�����(��I����*���$�QЌ3h��^(1�wHpF�Wpw�{W���)gq���;YEb����v
���X�z����d�Ƿm�6X����+.U���"�l$���:�L;�7��Zǎ�{���s.�k�Y�νu?~i9:0�����q��!A����q�#���W�+����CاWv��ycO�L~;�S�<:�諾;w��a�ϬJ��*fй�7ޜx�<���6Z���������+���T��+,��U��7z��ٻ���~!f?�������/�q`�u`��@��4������'-v����Z��^Z��԰v���'49�Ԥ���mشi����>�7�̈́�XZF�;���{��p�W��+�ݸ}fa٬N�Z,��u�6��ˊA��G���PD�K��J���R'l2"?��L\�����xb��[�49�3 �3��p ���Ë̀^�����o�iX"���'}���6u3�>�e�d��n�X�ҾM��¼ʳʅT��.��~�����@d���J�����./�(hzu�RA^���฼�'wj��
�����?M;�4�`�+=����~w�ϙ�ԛ�֩�,�w#���Z�/8�a�3>�P���V����?1خV�*�����~(�%P���V��<��_�Ӣ��w3�������qy���+��Ho({yzk�ҫW?v*bg�'���L�������u�g�׭��x�Ri�����U��O�?�p[��+�sx&^��Ppp۶�����V�>��Le���+Jh0�X���"h��B��:���::d	K������zI�Fޟ/u�w�$I�� �Y�}L���\�׭��o�W#|L��yu�ss��jH���#@muBo\vs�w�@6"��c���@�ie �$yK־�h��Գ�}�����ߢ�׮��-��͘9o���ɪ��7VU.ې�����pz��k_��>�'M��3����.�/x����Q����.+L��U�rU����[��:��B|���Ձ��
���B�v�*���ݕ�6�����>�ZP�/��O�sm��9f����&�#��lX���7�)l��/�.W��%j�?�]�~�:�ܥ�ՅlE��VY�������;���o�����zA�'�Q�!�v�!!'lme���o𻌔��Xi/!s����k�����S�Ol�.�+k;>}[��m/�d3�4�� ���F�-�Y�ub��Er�ߩk�/x�^�ͨ�MS���[�1���x�v���%Od3�V�G��I52HXc�6�1������Ĵ����_�%b�m�F�`HB��`�)P�`IbN��h����Ԉ�!i�F�}J��Or2(�x��$���W�x���>��E���2�/�S(�OZ����MqF�3a�Ĝٰ/#�'ѓ��8�� �w	rĿ���\(j���������]�"u���������#�J����T�W��������@$���-E����<"����F�{��i�^�u���Fp���u������i���|~��u�P|���,X��zW��O�4|6k���H��xɜ�����벗<�߯~�}�����O��0k���>�*��i���i=�ئU�	u�#�pҚ�%xRD0x�iѱ�6yӻ�>|�X�K��ۏ�:|�Α'kkOf��Ыsg���"��s��X!}yW}O=o l`�,U�Y'��\�U����I���9��繷& p�`KowsH@�{+AMg��#��3641�ı�au�za��x���Ӥpu�:R��Q�)
A��1���[�-��_�Xr�����$�R[ۨ�F;��$�ڐNV5���������k=?�g��	u���q���c�=�b�G�A7hq�8����;㐝}�\�U
�=�o�m��i��v������τz���{�qI�r���ԋ7!���˚s��R�xg�zM��V�~���'vN8y��A9���7�6W�b��^������;�^���m4��e!O�TF!MV��SP'?;�kQR��F�{<C�o�~�'p?�m���;w���,?��t��7&!H�G����Y��k^D���;�B}�tId���y3`�	-��`�U(%FL�!8ƨ��w���C2�27�(�E34-��E�BK�|�h�=���f��Ik�`tj�}hk��S�LC��z�~��������H!�o i�zظ݃FBvM`�w;��ݨ�x�r�~W�c�w�����OT�����P�VNUn��k��Fi�-Gz���ڷ�l??���ʡM�-ٴqɒ���|�SC�ݟ��@w'�6�7��j����	�Lu���%x�:O�Q`���~G��:��D\�����ND1��������z���*w�z�U�w�������VA!m��v�T�Ft�yL}�5�A�M��Q���@\@��#�QA
5)�,�o��ɽ�1�K:@^B�{c���/L���z�>��Se��m�Y�\�������#��w��鬼 �����ݺ}��lV�T�o����������l�QP;���]xn���:�S�	C
���n�]�r�_����1"ǣ�\����G����N`8�z��N���By���Sm�.��0���R~N?����?���))Z^��� 6��0Td�kc1��)耏R���r�}e�#}\��u5ʦX����;�$R{�^{�N�=�s���Mk��KD@D`5��դ�X�ջ�u�O�ou�'ue��ы��F�@"��%�����\@�x��36��o���k��t��~׎?66�PƊ�B,���%9%��0{����:�~��=k:vLM�\����!{��P����ɉV�9Uzmt;��E_��1��$�m��o��ڡVx�;Oa�YЋE�/��!�ԃ�_�h���-m�:��ܳ�o���1����t��K�\&�S3 �}��S=9*m%��	�'d�­mL+\���
�cޕ�\�t�o�&$Ƿ=��O�z��	�vI��HU��Oq0fOlJJX���5qCt��]q_�	�o�з���8����=��2�� �̚\$�٦�ճҰ��~��fH&��=��p�p�7��<��h��x:��&lc�;7�=��Iu[�hъ�-�Ƞ׭L��^����:t���K�^�ӓr�z�!�Wa8m���`����[�������3;y�(���Y���GMT׸1����ؽ./��@��ff,��룻3�����^Ɩ[�TÞ[�h���#�~�o��Ax�p+l�V��[_ݻ��|�#ȭ�	R3c�ဌ+ы��q#i�@2)��9{�<�RY�(�"y��iN����W ?������������k���'&g���V'����x�:�y�>;�����׶��X��۩�ϻҍ������t�KG_$��C�aku����VsV�%���ki߭<ISl@�ۺW:f��%�V/�����?��M��������~[[�>���{����o������vm��n�k�3~��
6਑c����_[!�P���+�jW�1�{����8�����+���ϳ[��U#V{D�`mߘ���55�w���Ur�a(9P���?5,�=�M����m��9!�X}����":.��&:cYJDÌ�+(�~���Z���1р�QF�c\X_��/�M�X�z5�!�np��a����������$= Q<�9щ��?�%�"� �y�[CH/nd���������W����l�x��{�-��p@��֎>nNLA��ʊ���B��=�kV���a���>�-����6qA�;���҇�uO��jc;�wt}���wh��_�#^� |/��`R��D"�"�����3�w`��m��~��<:�͓���y�yN��W{�n��g���6�ۮn���j� ���޾�AYMZ�ɶ���K�w�OylG��	�^y% k`b�9$�z�a��]٬�7�%�o��+�8����F�Y������k��߰6q�0~���4D��ȥ�JTi�����[,��z�G��\�ፇ�Y�W�fM��5kV����7�ޥW/t��O/}ty�����}>��0�P���Gԑ,�屹��]cl>�����C\,"�î��������f�ش7�������nķ�h{ؒ�gd��Q�)�[زΌ�?�ۘ��
�~�䎒A�3E�����qR`d�0_�Y:q�7�k����݂,���"ps��Y� ��=��s��ǓX�ʚtӚ-xlf®@���S{�a]>9��!��鴹��8r	t#=Q��*���z���͘�~>"��B+�1���O�;�>�f{-�Ln+�&(�g`\'-L6K5��|��h-��tS�6[&��cbN�����isf�{}貕u��2�p���?�<�������'҆rm�y��CAAGz��=�;q�_;��=�� {���}w���dp��;>n8`48;0��k���N�Z��?�k��w������W����;��#��_�P={������z�Җ�o�k������Pp8�k���Z��k� 8k.И"���y����o���էw��;��qW#3~޺#3�KM���c!��d�c����HkL$~����~k��8}�d���X�S��&�~��W����n�PБ�Ӗ+?��1���U=�����8�UK��x�Nw�\�$-��g��u��ZVd֚2�_$0�΂έa�����Q1(N�Έ3�I�I0�q&���Z�|x-��C�}��8-�9aY����T<C��|��F/c�i�F��	�s���x��\�C��p�Z|w��Ć�5�-u B|ԧ���� ��^=P�5Υ��y�����ν�=���������ŭ���K���ru�TN��o�nvs�.�G�k\+~H�>�Vѯ��/�*�o�mZ_�6���������k�u	qq�����1����r�BW�}`҇s
yI�������>1n��|'��'p^�Q�^TRҦ�,�~-�x� ����	�I��(F��ku��j9��;�}��C��l>����ɛx�0J��Ԣً��f����\�|�x�*��=�{H6"�[!+Բ����ԩ<9ib?�B6���+�L�Jݫ�)tnMʹ�Y���5����=n�2Ɯ���I#n���X�̊u50PHV�M�y9)�XN�
l�nq�.qނ,AU#QjE����U�������`�S���I������4�!�e"����G�|��S�6Jv��7}�c]�B���gw%�̓.�m�t�Yy�\/�+�D�U�A���$���Z��N�N�N5FdL7�1�qu�(J���4Դ�t�t���e��iW��[���1�ʣ�<*�ʣ�<*�ʣ�<*�ʣ�<*�ʣ�<*����e���G�Q��gAyc�ƿ3���Ff���1T��Wa���C[B&T��e���m��+��3j�^��.Nk�z���~�0s��#�����9Hodp���C?shK��y�ޖQ;�,�m@��s��3�r~Yo��
19�mW����������-��:["#"zX&Ͱ�䗗���d�Z���,��T>�̒�S�S:5';��3%sd�%+/�hrN�%�4ǒ_d)��T��e�..��/��I�,*�/.*�).~jdNiY~q�%2�G�9̟�s��`�rX>���$*<<��V��W�f���N�	+�)���T~x~Qv��������������x1�S�9j��ҩ,'�2)��xZ�0��=�hl�4gZ4̍3v���񿗭����@���43;�0��)KqnK,FcJNia~�,���)́�&�f��d�ZrK�y���B-�Ŗ̢�PL(�T�M�U��h>�</GWDfVVqa	��� {�&iK�@!��΀,ےYVV���	��*
s��3�9=�� �N��`I+�-�2�,()�))-ή��h���I�9��fBAKYٜ�i��y��@La��_���V��x�N��0Gp-�[��F(_3���R�z���@��~��9q����\�XhZ^q��r+J�`�11��RVj)��4%'���h2. ��ee�s>ʢ��tx�9�xj��@�"A@���ʴ^���&ОY��2��I9�Ԁ0��f|�]�Z
�Ksʶ�|FINn&,���ia����8;?7�ZfA9�4 ifv��\���R��� �T,��S�?�H�1�`FI^��-43���vz�Z��Y\�&��-����4a�
fX�:�T�ÿ}I��2.L������hL+.�.�6�b _����]7P���G'���c� =p&��7�3��ƒYR.�9� �?���-��Yn��,�9E���5Yx��B�FW`��q�k�-+.��-T��i)���>�$3�����bQqc�����l)Z@bNA.'jH�%>9)ݒ��>*:5Β�fIIM�k	�N���P˨��!�#�-0"5:)}�%9��4�2,!)6������fIN�$OIL�����A�#b�[b`^Rr�%1axB: MOSuT	qi���AC�6:&!1!}t�%>!=���і����A#�S-)#RS��� G,�MJH�O�U���hPr��Ԅ�C�CaR:t�Z�S�c�G��&˩1$����|rڐ��DKLBzZzj\�p>�KgpR�p.�I���	�I��8`%:&1N�X��0<�=<zp\Z�"|��N�8���qIq�щ�����A	�rLH��.F��A���A�IiqO��g_2$N,DÿA�2�~���'��7�2*!-.�����I�OMr�>a�qȓ+/I����=h0������N�i��Ƃu�M��))維;�E(��g��Z-�	.���D�<K�<Z�kr.�%��ᗇ�n؍��=5�`%��<�L�/��`a���e�b0�q����V�Hfs��o�%��0eZi~9Kf����Է�R}�j�_�%��9e%�S�O�)�cK�~&(�/�,�Pg]�/�<�C�-��l`r�0��d��@�(MFy�YP'��:�5E@��I0b`L9$��0:e�B
�	�Ƈ���)�bA�����]\s`�T��0҈b�50�D0"�f��b����,�1� o>����bX7S<k�'M`��è"�1P��S�_���H����l�}�}nsܹ�W�\�sX�E�?����
��`\1\K�׳𹥂�0��s��4��)��>w:<-�%З(����x�����A��ge�s���a��BC�k�&�
�a+kr΄�#�ژQ��������wح�7x�ץh�3�V�T���b��ߢ�s�"�
lM����rt�&�U��=f<��iN�j��5�t
����+��W���V��Kڎ�\P��#2�q)ѱ�1����l�k+��J��2�/X���?Ȟm�?���*�r��.�\h�vܩ�Ʀxt����/hv�Wl�	�)X�T:����[�O��S���B��KY@Y����d���<!�u��>G���K�Y�Fm��a��vx�P�Ӯ�&�-�١��Gh#��"JYf�4���T�k�׹�KN���Ѣ�[X]Gӄ<
�
vo��H�0�a�l����%1Fd	|�G;.У�]CYb�lAq�Ni���t}V&`,��I���IF�����P�l��WJ�Yϙ��&5�m��i��"y��X�H]����h���!��Q��k&�_��e2���B�}����^�G=�G���4�A�Vg߿�*��* K��g�([P��U� �����.\ָ�=�f
��l׾FK���&O�1.���e
=��_���z-��0Cu��y���K��#�+l���S�h�v�i�����.���	������싁�|�����w�@k�|'��>3I�}���?�51��?Db<'+��>����e�Ț�8�Q�Ϳ�1y"�[ĵL�1GX�/ۋ���b8Z�g���
��|%���[�-�Ӿg7y�ݣxQИ���3�c,��ɺƴ}�Hȶe���E��e�&�>R������:�(	��:�p��FA>�*���@>�
OF���B/��	(�q�9�d4B��p��GC�m��n�O\|n����b���m�������c&�/���=�lT[/I|9�E�.h�(M���U�S� V�S6�R��i���D�k�X?^����)�2�9�A@Q���#��"��!N�#V�6I��5^��&4��?�?Z���?]P�WJ�G�
9?�b>_u���(Kֵ��MX�tYjtp��l\9M��"�O��t��h�o�k�����F;!��rH+Ĉg\�\���#S�2Hȋ�S+V�I{('vl͵�0밯0X�'$�(F���`|Bc�f�	��A�l5���k6�� �A�G��'`�8ݦ���s�y���M�:� �&�'��Ԩ�daeJe���81*Z�:�Q
���딏p�0�G����HYs����>����}������S��(��ƫŮ8�ײ�yG��x�k�s;f�MY�c���b�c&�E��bla�qM�Z|����3�c����~J�r���מ}h�[;9f��"O�r��ƬD�?�3�i�iӞ�����^�XW�B����_f�l��V�i����X"�{m�i�]�g&��
},���T\��T�[:���[�/�.Aڙ*_H��a:�Rd?�5ɄK@{V�B�M�ǱE��y(��dʳu�k����F��ď�����6�����A�Pw�����%��d#�6�M�~������Fv@�U��"{�����_��>H�A�-r
�o���}����6a6�-A�-e�C�<;��hȾ����_",�e�8_3�Aش��:"����!�;r8�F��Crl|b:
�,͜�"�f���'��<�R
2�-h\Afyv���M�f��"BBF��Rc����+�l�{=�!!m��&`��Ó&�6��z�K�P�4b��G��"`��=�*|
E��O�ߨ�`
P�H\���	��F~(D|{��`Z�2���k���逃_�6��Mڽ�l����&E��mjx{�=���X�]�v����$�II�5>�-p��	�<AY�s#`4��,%�C���F�Y����e��a�����Co��dS�$Q��8`2 ��V\ �WO_�~�c:��{"l��e��+c�ۖ��ƞ�t[�f��&B���W��m���وn�Hp��2jɡ��#T�)E ��:|���u�6��U���7iGI'Fz�(b%�$���2�d�)��L%�ɳ����:��j���"�H9Bj�Yr�|D����ur��!�)�25Q�C�hڅF�޴?��ChM�c�D�Kh)�N���r������V�����Az�������9�F����]Z�30W���0a�,��e��X6����l���X+g3A�Y%{�m`/�ml'�����8;��c�e���ձ��S%&%��-���NR��S���R��(�J�x)[�"�HS��ҳ�Ri��N�$UKۥ]�>�F:"�Jg���G��+�tS�#ݗ�,�&�C����r9B�-��c�!r��.��'ʹr�\*O������5�zy��U�!����c�)��������|M�V�%ߕ��W�Si�X�%T�T�*�+��P%E��]g�g7\{�Hf�m��[a�3Rn˰C\�p��V�y��^h�����o�B�:�!`�����z�E����m% l����m��6Q�������l���Tg7Ґ�r���:q��Ī��P��@'��p��t��T��!��c�x� �_s9zٸ��8�6��
���� ��p�.=V�E�f��(cD�D��k{��f��=	�=�j#{
8L�<�!Pr��lV�w�ӑ�/l}.P�$`��d�x��#E�����_h�3C@��o�+�_#������b|mS?��pH
�N	��;�-����l;�5�m0�ko�HV�r�	xvN�' �	�c�'�Yh_X�^���l'`�Z)(�0�K�@�Ca�`��4f7�����t[9@԰���Ԃ��X���Y�l���4�~(ć��T6�����pXȁK8C5���XH	�SA�I�i���tՓ�����O,��薀�8��s��y��+b�̆����@�x����۶�~v�q���lОb��窾6��/Ǡ��(�0�l{BP�w���'��_U3�%b<`��.���6/�ǎb���Nr��m���T�`1<��Gs��i�����0�9n?�p-�(u��BA��h�ŜXn�����)�L��`!����G�\�(6
���"�b��@�.�QS�)�:���2�c���4S�i�n�7�D3M� ����}��٥3����%}����z.�ޯ�2�e��J�=c�=/*w���[FW�~�1W�����q�g��i�e� S�#2�g���-����pҾ/�Od_��#�1�B��u$j��='=Г�����V �T���§�9�����o�-|�Bĕx�6�BBH(�$}��$�%)d$G&�<RD��L2�,&��y���g��p:9@��py�\$���RGn�{D����z�v4�v�a�'��VOi*͠�i6�BK�T:�>K��Ut�D��v���5���g�y��B����Mz��g����<��cX�z��,�aI,��aY.+`�l:X�B���a��f���`��~v�c��9���}ή�o�-v��KD2H����F�H!R�)���b��R�4R'M��"�\�)͓K�����%i��S�+�Kǥ��{�E���T'ݖ�I��d�l���vr��I�{�Q�U���T9C/g�S�y�<[~V^*���ɛ�jy��K�'��G�Z��|^�H�"%_�o�w��
Rd��J�����K��s���[����U�M/����㑟1�1i��g|>&�́�Yxld��+��V
�qO��uڨN��#�ԉ���X:�z�S�Y���$ȑ��VP�G�c<���I9��g�/��	�f�]`	�;��C2�Ӊ�P�o>�yQ����"��;��F	#�D����D�J� ��<y��`��1��t�W<
8L��'9�k$�K_v�KU��A�[�.�Zc�$��_p��$C��	�]�������Y�C�)�X��O��p!CN�NvTH�_ $����w%��
�_Vr	��/o�C����!�m�h��! בg�'�A�{�ՙ<o�0�RJ�mnQx��H;�-$T�{\��˭K��Sd�!�r0�6����6+m�z8��5�jE��ee�f�'X�l'
K�4_�֎˅�O�6��0�-S�yL�l��p��s��~"���1c��8�%(�<�$�'��Ƴ�������l����G�����?ГªAh��s��w&�?�gh%�@��i���9��N':��ɥ�,t������O�"�ׄ?���E��*:�����zǀk�D�p~��_��ΓE?����=����K�\Hx<��&�����b<�B������o~�$}=F�Sh���l�$g������rmN�<J�0��9_���Kh*� ����T���K�Dҙ��#��Mʳ��[�c�3���Yx;�L�����O=�i�&pj1�����o=�}�[^�x���0���a�A&C���e'�WP��t�L��g�D>S`z��
M���<�L �̥#�3��|��g��߱�;u0��9uA&�L|��@��қ�'1dI"�d�HrI)%��3d!YN֐�d3�Jv��d?�HN�s��	��\#ߒ[�.����+��m����PI���i,JS�H:�N�y���әt]L+��t}�n�;�^z����i��H/�/�7��ަ���323�f�X ���XOŬ,�%�T��Ƴl6���� �g�R���c�X5��v�}��a��,;�>bW�W�:�����d�$yH>���A�"EH���R�4DJ�ҥ1�D)W*�J���3�Bi��FZ/m��J;���~�tL:%��>�>�>��I�J���R�Ld��*{�md�"�ʑr_�q9V*��#�q�$9O.����<y�\)?/o�_���;����|\>-�'_�/�_���u�m���*L1*f�[i�*��0���X�x%QIU2��J�2E)Q�B���TY��S6)��ve��O�Q�(��Y��rE�J���T�(�� L��������a�m�o�11$ �X�l�5�tў)�ɢ��C���Hѣ����ĘkMcp��v�U�t�c�O9��whOuĠ��#뾡��c���V�Ǵ��s�V��7����6m�#G�5>��H�2�qO��~�R}��*�R�/�Ru��2�i{����v����38�=�MM���m���j��c�?����h��L��m�rtJڬ_K�=�͟j���9zӃ���B-Jh��h9�������_����4�t�Ѣh���l������+������)���6b��d¦����6���-D���r�A�H¿[ٟ"�9˓�z-A=�r�E�M���v�4
D�Q.�E'Q1:�it���+�k��w�=̹�~@/���'T��z�ٰ�6c'�
m�޸5ڃ�`�����8�@o���)�6�����#����"�ί8����ίb��y/fί9�ǒ�E�KXq���*����=�����\���B�'��7�g�$%O)Rʕ��<e�R�<�lP^R�);����r\9���\T.+_(�(u�m垢��h0����N�0COC��j�7$R��l�C�a�a��Y�R����3l2T�v�jG�����W_����>������޻�~�h�jԤ�PeǠ1�C%�J)*~`RBiB�Zk-5�j�!�c�!F���X�fcm��q��8�Rk���c���O��x���a~{��ww�=���%\H�b�^!���PJ(-4844�����X(Q���(A�!*Cաe��x�,�Q�X�h@lB4#�#v�v��^B�hm�������PG�"�0�h�aa��é�a��q��ng�a��0�p�9����Qwm.\�(G`_^�X��A�A�C�#M�-�Dkxwx/ #�!N"�����x���ʘD�eSW�'����C8b�#c��r�<M.����C,D�� ���K+dԊ���B�7 6"6#�"v �����(�$��q��|F>'_@~�1�s��N�LD�����a(�ׁQ0Ӊ�ɀz�#j�ϔ�*���JX�� u�;�;1�E�P���CpN�i8����ԝ��SPw���J�����	��0%]A�)�݄)Y�$�L���|jO����r:��S+�9��~G�)�z�QiRPg
�LiE�F��ԛ�zSPo
�MiC�+�9�]��SQw*��*jOE�;u���Tԝ��SG�c��j���NS�"u��P�P�Q��+�U�Z�NݠnT7�[����u���zD=��RϨ���e�i�4�L-IK�Ҵ��P-C���&j��)Z�V���J�2�R�֖i+��Z��^k�6i��vm��K�@ۯҎj'���Y�C��]�%=AWu[O�S���z�>B�Գ�Iz�>U��g�s�R�\�����}��N���&}�ޢ�������~L?�����y��~�aC7\����h1�#�1�x#��5�F�1�XhT�K��*c�Qgl06�����}c�����8b7Ng�s����^&���d��i�`s��a�2ǚ���3�,4g�%f�YiV��̕�j��\o6���fs����e~`�7�G��i��a^4�X��`��m%[�� �^+�aeZY�$+ǚj�[3��V�UnUY���V���Zg�[�V���j�Z���^�u�:f��ڬv�uɺj�ۮ���o������{��͘����(@����6z���k����6��6����k����6z���k����6z����k�����q���3�s�b��AKuЋ�b�t��'��u2�Q�Xg�3ٙ��9��l��)s*�jg���Y��:�g���lwv:�����!�s�9�u:���Wr\յ�d�n*b�{���p3�,w���Nu���\��-w����r��]�s��F���ⶸ��nw�{�=�sO�mn�{޽�^M&��D7�ob�āި�����o#�͊2�{�*��칞x�7� ^�e���t���p;卵n����G�����s#��(y�+��r���_�ܫ7�xzt��^�Ѽ�{�A���bݝ���j�����گ��~-w����{�|6��w��3�[Z�o�����swҌX��U����Z�kz����i'���x��u�Z|���o^��y+����|�k[�ߣ}�h�%��)��/���=��u����ݷ�m�ȣ�s'��i�:�k�K~K��<��+�O&y��oD��21{�Xu�l`*���WW@< E����ѣXwF�X�[��D���<�3��=�5�k�왮m'y{�<�<o/�V��u���-�����m=��H>(�6��<OD=O�l��9�Z�.*Oq����(OYT�w��K��IueF��E�/R�R⥱f#$_@�, y��<��dE=��g�oU�x'�֑��o�omW�b�z@׳��gS���t�����fh�g�U>#΢���ETע(^Iy*��$o��'|��`���x_�}��_[��sH�r���&�M��r���S= �I<��'�js,}uنN���<�K+�$=M�E�c��u:���w�u����Y��Oz6҃�}s%�' �x.�q��/ ^@��x���WK�o+��[��M|4��ħ/&^�e9~>���}������;?��e:I�����"��I>���ӛEyf/$^����z�1����xq���#��k����x1��)��TN?*�����z��'�4�F���Lbn[	Xǆ�:��=B_��=l/[���VI��_a���U~y�$����7� )���I.9�(>Rʔ��R�4�ϡ��%�������xE���Z^x5��W�%�%��q������-�[��v����O���7�����7⟋�o�_���__�7�j���ro�ߑ��-�Z��V���O���ҏ��}�S��x-�"�zKoI�,����S\�=�u?��_�*��q�X%<����2���@��$D
���·"pN�G!��$�MF�=yb_�$^B�X��Z��A�D�=N���A�B4��K���]���~ZI�\��:�u�F�Et�;띾�Գ�����ֲ��>���S[�ڊ�����|C���3	�:�>�X��嬆�A/�g���ma-��h/;��c�$kc��G��U�a�s�����@>��#�>�g�\>��">�/�������Z^�7��|3�����ž��\���t���c_��`,�r	�ۂ`"�P��KF���a���E��&!r��*1���R<�=}U���'v�a�ڧb���t�ׂH;�}���j_Zx+�a����E�>�c?��L�����9��>K)���y3�3.g�@�^��y#RӋ��W�����g�CNIe����t٘R\hŅ�Q\hŅΦ��<��Mq�y�Ge�~��c�H\I�~FZ!����f�̙3�/dYE%�sؤ�ť�YNqiq9����,�d���s�Ν?��������T��G���Gj��4�z+���.N��x�2Kb�χe#�61k:7R�4�!����ŞN�b}�;�����X���q�W>�+t�ѫ$b*z�%Z�E����x�F��EZ&�l��;���;�a/3I���d/2�-鷘�Nڃ��.I�P��"l�K{9�'�	E���{�~�K�m	O�k"�d!�hx�q�0<��7�[�|��,���$̇����x��O�g�x^�_���*�o�[����o���������ā$�#�z�W�._���i��h�e8��M�+w)���8��v7L�G�q�6|�3a,����#�1�~���Kx	^����ޑ?�?��&�C�T��X�5���kp�x��� ���`zda���[/"���v�؎,)������c<dC.L�<(�P
ePUPKa9��U�j��6� h�/���6��|Q>a�*��UH�������Y����cha<L��&a�/Q�'r��=�̆�x�!؊�h؂�7μGg�љw���R�ɣ(�Fī���Sd�¶�$�	o�a���e�rŲ�L�D~��������݃t�8H��&�O
endstream
endobj
20 0 obj
<<
/Filter /FlateDecode
/Length 458
>>
stream
H�\�ݎ�0�_e.�+��D����H�菚�pR�� �\��k|��H���4����ƅ�q�O~������#����:���_������T%��y_��.��T�L��%>��m���U�������ޜ�>=������І�I/���ߺ��*�^�CZ��k������=ɬE������.\=�7�iߦ�&��֍��|�w1��z��M�mޠ�g�-T��j��P�.P���P"4J���P
� ��A B� @�`�V0 * �
��T�Q0H@�� 4�% ���iͣӆG�a��Ў�Q"���>�t�#0�G`J�(1�5-��Z��‶D���ḶD��l� ��-o��8��C��,�3@��9H��m: \i%�W�����.�O��u��y����cм)��\gr�cߘ�yu��  �<L
endstream
endobj
25 0 obj
<<
/Filter /FlateDecode
/Length 14523
/Length1 34888
/Type /Stream
>>
stream
x��}|Tյ��g�s&���+�+�$IHe��< Ɍ3^��O�(-�"���H_�����km�^h����z-�j��49���>g&���m��������^g���^{���^{�9�㌱� *sW�>s�s�6g;`vaQ�wzMc��ͮ(���s�|����^9�ja�g�	3v�P�˫��ޑ��m���h����ퟶ��a������[r=V��(Ɔ�B���-WM�����3h�`�;�g$�0�FC���O,��r1�?��u{�L�+�%�&5����ml	����?��1�}?o�չ��{�ǌe����Z�k��ǴZ�ߌ�Vw���'N����q[��C�M�r��N����_�����򝑺R�8���/ѯL��6(���gG��\�[���6�m�J���������g��JJ��0�i6B�N$�<� R�X4�W��t��׾���*~�ꕞ��t�]U��~���� 4�:V�y����a=�L�;-����~W�
k��2��'}/̆�O�u|"[�
�J>�?îbW��X�m`�l+����61�Y�L��t���v�[�~v���z����>[�ְel�M赔�dS1l���@e�����mGߥhw�բ�V�C��D�uK��|�^V����t�<̿b�a|��.���� #U��������|����O�=�3l�L��{gb�b��ډI"iM�,��R���w�D��j�Z)C$����J�!�t�zE4���V�!���b���`��^�>��1#[������ÿe� ��Ho�l1Bm4B��07�vy݄�ؼs�+!��2}� /�z��C��ẝ�fc 3I�����3��sk��̂5r>zI˨�mdH.U�6��d��q����Xoɏϲr�	���VXqP^����� ��I_$���_�%mXZ?�Q�*�}����7��gϚ�����K�ѕ��(mN=ZG+m}˶j�d��%�?h�a}�g����@f=LE~��"m����+gt�=��q��V�®a;��> �Jv'r���M)��-�A��XqO���H�,��+f��t��aY�\���/��^��N���fȿ�5�?��mH�!� ��[�6�M@��<�M�<� ��"%�8��4?��.i��>g�+�|e>��=HT��7�hWʏq��4���p>�s��Il;���^�s�!�A=�`�R>t�����?�]�:/C��7y����/���
^��e�~��j�)	��2q&�J���`>�9�Ϣ�>�����-����i8	r��١�+�!x��7&�Ƽ�\g>^h&��������y8Xz]��3]k�C�?�a)��`Y��DV���l-��K��;�V���k%J�\�y,���aE,O��E�c~��2͡,s��y"[\�����`1�y��@�~/���w��E���J�~=vH�Ǟ���������C�@�(�Aj�n�(*��8���yYR*Z_<cU��|�x�]�։��r�C�c��%w{a��E7����� ��M�4��R���#m�7�!Й��c��G�f,Jt큑6`,����C�m{���2��x^)q�Iɕ�e������1�N�.�؆̱~�� �"�$?$���2��06mi������Fy%�1�Ay�,s.�<`�c��6�1�+����x��������ȳ!T`�|� -�c_��+ka�[�վc4��}܁�n���A�}����6�X�>�l���b�LG� �(_��d����=�0+Ef�h�0r;
��}~iFx�������s؜�{��r�alv�ð]�8�}��!�B��Ӊ.�~�7C[31��AK��C�D~�mè�c�5j�s;��t#�gb�7��w���V�s6�^�&V�nR5�D�W�<hY�<�'��J�U�;@{;��x����'��_�;�x��R#���C����Q��.�eMO�����>X���Q-���K-����
v<��3�(kGF�3�4��ټi��+���I]f�\hj ݎD��*���"���f�>|>h�#g�n*�����A�B��a�|�l)��ᡇ��\x�\��!G$���V�2��8�ɾ@끠6 ��~6|{xȔk�b�H�DU�sldu+RFT��Hv��o�k֊�"�[,�R�11�̴N�R��TL��h�|�T��T����!�B���8��g�!����ce��M(���46�S�ي�<�[J
�ӱ��N�*sb�:�	��=�]�p��S�_l���c��*���|�|�}{�����a��U%����1���q����<s��0&��/C���1�:NcvI�����t</�%���Q��ef�ys��x%n~�%�R���}��� ˷�3�S�_�b��/������K�N�?��`��eA�	�FZ�#���	t��v$�Ʊ��ߚ�fڏ��+ʏ9�EA�z����/�kat�-�%����0��v�v�]��`S�6��_�d�_.�{�C83���}8�e!�n�x�b_a����IҠt�uS��5�#q�Ċ��Y�}p�A�/�~ϰg���8	g �ȕ��lF������z��ir�ɕ�ϵ����3b����1Y��ӸA��T�f4���?`�tVSW-G�4���%�'���T�5=�j���}5d#Z*�B��v҆�����ȱ� �ʖ׮T�5���Q�@���e���A���Yg]�v5�*����%\"�à�=��#v�m������i��zldg��������-(�,�ƞ�{���h/��i�wNʍΔ�"�Ⱦ:�CM��]h}]�����L�V(+i�e��;��Q��!�iX?��c���Jp�#v+���.�x;�\�9��t��D�	az���3�>���S��/���Ֆf����7	+e�=���(��!���sx����ا�m���L�C�=,Ng��}N*��y���W%� ��6翏���+E���kq]��F�=�ܤ������F�A�FI��NJ��o�'�b����|��I�Cb�����p���KU�����T�ԥ��U�_ß.cӇ�t�5'"/�����<��h���v�w*|���&�2t��ho!/=1�����V��]�x��^�G� ���Ѫ�{�]�����wYo��CXS��7�'&��v)�.�����%��f�g�qֺ�V���q�i`��FFqK.|��Kp�	 [	�.�ic2���8	���)�pf����r�͈I9v�3�vDt�qJ؄S/�Us!�(�GA������ZN�p��]�����<��	k������T��v-�iA���G���6�e�� �I�0���8w���	��Pp��>����ag�ũ���L���`G+���|��,�+h)̎�n ;�%�[�z��g��W�^d/�_"�e�y)$��U�� �����)�r@/�D�+��h���Q�6��(����,�a�"�.X�:��H�8��x
�k���A����KF���K�w�K@ܝ�VoG� �
yV���]�o�q�vVT��8���`*B�J&�g��"��o��O e3�rc���®�eQ���{���.��ӾB>~�+N�+(�,J~���W���}H'�oI�,�0]�8�?R~B'@܍�1&�ӑq�Ǚ��&��������?��a�;�t���z�w����ɷ}5?4�ߋ\���ᷣ�9�Zұ�Q� ړ�8X���>��?��y�x��B��<������'0cV��䰭�����K�+�#|��C�<��.Nّh�Hr��py�p��a��I��#�qr����!dz�����(> X.��ƫ��P�k!}n!|B	��ʱ��D��Q�	�@�R�"����s�zE>���'V����)����,dz����;++�B.�3�A�G�\ng�٫���'!_ig�X<v&Z;/�^tRr��9�r���^����Sc��'K�U,i�e��0f�FH����W-; ������O��
��lW�aeX��pނ��K���v�Jv����=ֹ���5jm�am�a1,�:l��_W����y5��O�T�VWU�"�|Q���Ak��d�aW]���ۆL�-�;m;�l�3œO�'�?=+~rVy|�v�I��l�X�xt�x$W<�������Z%�{�Mq�_{hΊ�!�?�E�o��O��[�=�E<�Q���,m��/O�Q��k��sŞ��{gk��⾣�W���?���-~�/v� W۽J� W�2�=g�γ�����S��0�=]�e�m���)�4�Vo��u����T�4q��d��T�%Y|�>C�N����n~R���oY�m~Rlި�r�0���<��a�������������z�r���zi=�^���b�G\S%�ūs�z4X�+֥��@���5�Xm�P���!W�hS\�#���o�t����j����Z˓�e���4Lk^.���U��Jܬ|R4兇�F�i�\<�#�go�����po+Lq�G,�<U[f��S��\�dLOmI��I�YOm�)劅���rj�ɢ�)*�i��ł�dmA��H�(���ʶ��Qj�y��[�K��]��sΊ�gE�QT�K+� 
{�Y�"?Q\�+f��Kg$j��b�t�6#QLw�iS�hӶ��S���>b�Fu�SL�S'OJ�&O��ܤt1qB�6q��0>U��.Ƨ��Kҵ\��՗��qc��Ҵq�bl��*'C��N���c�*yy�j��$-;EdU�F�J�F'��G�Ӹ�'h�Ũ�|c�bu�<1"I�'���kYC�0\��C����bH����e���	�����k��?U�Od��a��h20WH������Bk#^��7E��K��x����M}���jz��3O��\�v�{�H�,z���Y�3W�$�j)gE2j�sERb���A$�.�F� ��p&iF�p&�����$�,	��aI��Z��'�(�{L��v������]��&2 �!XO��r�M�����?l���g χ�C�vv���N�2��]-~����}���2��CpFXf�Z�֨}�S��h�u&2��F(��5�j��q���/�d���V�Ee+�ր����b�}8)=���4�s|b�݈�� VSp}�'�V��������g|/�YPe���9�>{���^�v�=��k������h�~TOu�d>v�-�=�a�����]|;��+;���2]���e���N����`����g^E��^��Rv��"��������n%��^�^W.�Y	\����'2��ʿ;��|��:�z�8U(��ܮ6j{:X�<C=��c<N�UT6�������'O��+epʰ�)�U���onw$��2���O��	�`�pj��]�K>�@��r�qР$>	����x]MqՎ���Tpܗ���뻉�����&×�o�~�l�>�_r��\b��'O�L>�թq��KIf�s�����!�J�Ԟ�s'MV��\h�j>�g򜅻
K����я��2z�P~_���;�5���v3�_LZU`ULm�<q,��������O�S��6�GK���	F�O�L��6�@:����5�����pš��>d��g�[`3����_�_�;���[<����A�(�6ȿ�dUy����q����)��۟��Pذ5#}�s`�~��xT�S)=��L��s�2HlU�
5�')I"IU���<e���)�hJO�����/,|��|�<�/�c�*�yߊ����~N!O��tT���w� )l�8�:���������Q�A_N6$/E0?��k~���Iq,�H>q<��x.�)���\iJ�tP�3�G���G��p�loo�s+���ׁ�����LIR��:ć�������|��F{��c�v���F?�=���@PKЇ�	�؀������9�`q�y����z\^J�"�zWx���a����/ɪ��_.�|dk<���*����+���ʥ�eq��ߢlTr<��3������c�d������M|#�Ml��o����P�wO�^���w0�a�3q$��~���y��k��ai#���)S��ܟN�"���!���G���?�kb]�l=;Z=�Tn�{5��2�Rl���`Fz�~�pRk�@z���b�1<]*����S�8!9�2_��Ŕƫ�
46v\���*�7�j���_�O�0�l���j{|a*�:��\kn2�7��͘�M�ax��y3�z+}R���I�)=��ຆ�BM��4�7��/aS���_o�1�W*�?bhZ�A�iE������#�\m�k��K�M�/Q�/K2y�8a�����NM�3x�Tupf��I'N���wws�Æ��W_�*Pu�u�0�b~�{�q�4���(U�.|r��?�c�7�xQ����+xk��N��/���[2�;��m)��gyP]��l��pr��%�i�?����y�:�5��&�)́�+���?�g��{*c_��w�=x��
��wǎY�i)�:�B2�&�d��Tѯ11�1.�x+�>*KSrSҜ#�YΕ+ON4���S-?<1�<eJ2�OM�Te�>|�����y�>�_,�j�n�����+�l�(U;��]�'�t>��[n&�9zt2=Bk;X*����*�X�hL�ո3�G|s��.N+�����9=�Dޛ8�=�Ӝ�׍�4�w��{����F?�fFp����?3����]]qhE��r�ˌ��:�ƎS��P&�J��Lɶ����7#I�@��b��.���b��.���b��.���b��.���b��.���b��.���b�L�YOO����,򗘜%��*+Le~�,X�(^�)k�`!���^l�]�'�w�e'�����w�7�r"����$���c	��2g.�H���8�<�,ب(^�)k,�Ye�u��Љc����e'��|�.��e��ˉ����,�]���1�Q7ҕ;n�xW�:WAS(
x�-ٮ�ֺW~s���Z]�ޠ7����I(��t/js�5�[�A�;�u5���m��Mu.�����iS�n���Z}�_�g�7l�rs�O�P=U��j�O��Å�Dc(�6v���m9A_[��[�4xsZ���k�V5�mj�x����cK�꼭Ao��M<�\Qy\#�^�����[32��-$�IH����.�rTo	c.�IH��5��6rXt�n���X���w���P��4�vѺ��b����5��d��� 0���
�\��u.?�|�!��ڀQ��4�5z�p���Z�hNB���li�5"S�$s$�y\�`�W���x�`][��5�?�M����(;��|��5�y�H�I���<mu^I����j�B^�C�٘���6q��)��k���&{ j�T	�mA�'q�]-^)���`cv��4�X_��bк	���w��Y?):d�N����rn����@+�ʎ�+��v�jWz�B��t��$��|��&�#8-!�U�Z�j����"�@�Z}!LC��Ҭ�;-��s���kkl���]����.�_�{^�]�u~o��XLu�mq�#�->OS}��9�CD����R�/w |�5�r �7���*�hh^�oR'�Pw��G��`��,��X
s7��F��ᥓ"Xlm^�j�b�)�w~ɶT�2in"K���Z��<AWft-f�ؑ
W&-�L�6̎��VQm�<��}MQƼkCX5.�ߏ%�m�R�%?(w��Fw��������^0\��{\mp�_�]�J�%�f6���-��&��j&��i�w׭r7@0�E��������e(8-��m�'�����˪]U��Ջ�+�\%U����E%�E����*�gf��T�)_X�B�����%��bW~�׼���lWQMEeQU����U2�������Y�K�f�
Я���UZ2��D��eW�TIQ�_T9kn�JJK��d��K�ˈf1��*�+�Kf-,ͯtU,��(�*�B�-+)+��(E� �*�XRY2{Nu6:U���/,��_9/�8,�ȕ.�$\���hu���_Z�*(����,ʟOmI;���瓎��W����
� J~Ai��D�U�_2?�U�??vQU� ���S�avQYQe~i����hV	�ǒʢYղ%tM�Jvg��U-X�E����)�C@�|��%9��A\�S]^YeeqIUQ�+����X(�,�4��A2.�>i��l~i�w�u���,,�/�*b㜶����u^�l�^ܖ{������j-' �݊�k�d���%w��u..ڒ�m�K�֍��r���^x� ��9�5MA�ұ���}/�n�`�m�nF�`�ͮ*�!�M�&��3q�ۀ4���‽Uu��F����c�jZ�m^�����$'M���Zlѥ��B�">4�j��=�Z�+��b>��X�5�ֈ���F�:6�\6i<J�h�bhbA� ���d[�Z�>�|��\�2J+(Ｘz�g5�-X!J+AakC�:�u�J�l�B��@��/_�Ҍ�:�y�oZP]w:U�
Q��V��ĳ}=hA��'�悏�lr
����c����S/�-�B�&H�x�&����n��s�·k �{e߀�4G�D-��k��*�R*��~��W*%�Jμ�8f숞"�u��P]P�wZ�C��>�6R�����4�odK�n�by>�����G��?aîo���֢Kֻ嬶H���;�&^H�
I�ER�]�v����r5�QZ�=z$�zY덎fͰe{ْ/��U�������!{���UX��ٚ��I.��7Z�I���#���{s���ʌ��L9sn���|ա�ۖϲ�:Xe���5��뮚m;�s��k��s�S'���0J�䳓�� $m�^���1�~�l{-Ձ�6I���i��C�lʹH\�D��.Viq�&u�3;Tn������D�쯑#;*�X�\���,�M�V������h�����P7��h��G˷!�ꥇm�%�ƌ葐�Ȗ�6�ZP/$
E���q��%#3T'��H��lN���Ym������g蜃X_ԩ�s=�3!{5�����y}@l?���m�Tm�oGl�҆����O�ܑ\�ܷȫ��0��f��^z���ES�K:Y�E��&��#�x�^��X����:�<��"��b�Tܲ_D"���5F�e��#E|�[Z�e��1��'��2��8Os�9:��x��r>��yo���.����J�Z�Ѝ`�Qˌ����w�.3�FJ��3ϳ/fF��ރ�Gv��k��Ni�}�V�{_�m�z���j�6�Gc��콆Z���]�-=�7�#v�-�/�b��w�k���+-���Œ�|>�j��(2V_��W2���?�f�v��%���Ȋ��9��])��E�l�g���h�{����c}�T��	��b}TS�R]�����)�]5[�x�R���n\�e���z	��"d��|YC��r5.F�(�˗.�l��D{	0D�%��nڗ��-b5r�"�RjY)i���"���W!-�=�g3�F����B\��|ɋ�i5�v�D��l>�*A�]��%��-5E�(��6��RGD�h�G��q��/))��(��-�2�ޒ�Hr`̈́��,\+06��M���\�H�v�l)!�S(�Ө�$��ܞe*wRɱui�ᒯ$.�� �O/itI�����s���ۙ-)̏��B)_��C��@֑I��і�1�2K��8/�#�K�T�W����s>눌0[�W$5U*[WA�Eh_�X�X"e�e�֢iٽe�1ڝ%e��]�Q�l�ʗ��*��B��N)�ȷ��u�~�=���s].��\�,�k�H�ʗs]�B�\��m��XXd��Y嬫~#�(�����Vd�3X(���*��o�k��"�ku�c�k����ܱ�cgTf�N_	X^x�l�ҭ]'���֞�y才�ηsEN�VL��F��w[g����#�t+F�k��E#�5��sO�N�-�E�y/(ǵ$k�{t�eŗn-�h��h�B;T��_���(kd9dG&$_�ݖ�뻝��NU�4Y�I�9�~f�����)�̱�X�|֩Ҁ�]XK�Y�>�6�u�CI1�{���W�1�7d��V�-�|o�RXS�a��Y�����RX�-�+��Sى�=�Pޭ^͸z�z�f��Q~Y}�W�WQ~M}���0����S��73n<le��S��Ie�;�h�v�}�����j���kٸ�u�f6�!�]�*��>[���Bi��&,���*)� ��,�"���-+l�+���b�IX*���R�2Y���ل�yU%��=�d�$̒0�eU�*j�1���e)L����=ǒ3���l(�v�wU
�K�s�k+���������7Z�	{����5�~кO
�X`&3��\Y�A�C���n�=tϢ��2 ǡ5qj�1����H�^�	W�^�nTo�6Dv��܏Z� ��+e�-�b9{��XO�8	2-����{���>Ŭ?
χ/Ԇ�\���\~����Ť��3���t��+/���e�LJx��	::GBpn�
e�t���M����?��i~Va��JO%]�P�*��q�$e�R��Qʔje��B�W����V�V�Q�M�Sٮ�R�(��C�c����ϕ�W�7�w���ϔϕ��v��8�(RE?�Y"[�)b�(sE�X$��Z�(ZEH���b��&v��b�8 �#�)�x^�$N���{�cqR|)�SU�5YMS���5G��NS��b�T�Tk�+T��R������ǚ�C�[ݩޫ�S���G�c�q�WX�o�o��������Y�i�fh=�t-C����i��Z�6G+Ӫ���
�^k��Z�Z�F�6�Nm��Kۣ��i�iOhOk?�^�^�����>�>�>׾��uE���T���ҳ�l=W������z��H_���z�������-�6}��[߫��G���g������[�{���I�K��n:TG�#ّ���t�p�8&8�9�ŎRG���q���X��;V;���?>�LkH�3K��.3a�ʌp`Mxm��*���d���js:������L�0ө� ��7�wD����Iք�i��� ��$@#|0o��a�F8(�
FZ��G�����xV���_ґ��*�������t����(f��L�%:aZ�9z��l� �&IX�Ak貎I�m�8� S������!L����:��(���S��\*���{ ��w�2aJ$\,1�Z-'H8Ob��'5~w8�]D����YB_+a�f��n�+�v����c����Q���j9kh����;��� ;����1Gb&�X�q>�l�|>. ̖J�|/�������aO�e�f�?&���x��'������t<8՜����r�{���a�^�5h�%,1�4a��GT��({_I�d{�|A��"mLB��y`
�m,�/	��pC7����ar���煯t���D|���\��K�}���,	o�_Gm�[�c�!�-�`���*_��$?L¿u��������5x����R�yR�w�D����9��~T���,[Z��n Y��l@n�%�Ko��j�9ֿ��%~6iL�t�I:�m��  �,��x_��Ga�7��&_�
���2���&k�����g�Ae�9C���#^��&)&e�<OQǻ(?O�+s͙�?�-)���'�����.�q迨�LĘ.6�bd1�1��fAc�1��1f!�\k��8�>6Nb��+��ټt��f�N1����0[E�0u���0��vü���?��lⱏo�������M���y���Vz�*�:�Lf���~�~eI���o�0��-cv�g�Y��nШb�s�v@Sq	��4��ο�튢�)�J��Oq)YJ���LQf*��\�BY�,Sj�F�U	)땍���e��C٭�U(��#�Sʳ���K�	�-�=�c��rF1�*D�HD�!r�1M�bQ**E��Bx�J���5�z�Y�!�;Žb�8(G�1q\�J�,�o�ħ�8-ΪL�UC���Pu�:N���P�9j�Z�.UW��j�P��rnToS�T����=�~���������s��U�M��#�3�s�+�]S�8-QK��i.-K��r�)�L�P��Uh��eZ�֨�j!m��Q�Yۢm�vh�����vD{J{V{^{I;�����}��Ծ��h���	z����3�z�>A�����z�^���W�}���W������;�������>����~T?�������������O�g̡;GOG�#�1�1�1�1�1�Q���(sT;�:V8�͎�c��ZǍ��w:�;h�u�G;�z�;T��x�ve��,U����N�O���Km�>uU�J}���O�n����?V�s�\�S ?�; o��Wɳ����X:"%~D��i�ZA�4����c���)"E��U��AQ�jA�d���:�3�?{�R fI��!��:�V�n��@e��p�v_t�tq ?DPIV�sn�h_�K�8�$a���1�r	�IX �
	�P)�*U�C^&9���y'I+"o�Q�v�F'�j�Z�k���j8�(ӵ_�
�p���3�S� �:(�I�Q�]�I�8Q1�A�o��G�1�	�>|�J�^�÷��Q���C����U+�R$�s�:�?��x�����<���)P�.�ZD�i�uh���Y=1�B8{F��Ĝ&�#�Ս�q;�7�J�f��Ɗ��N���Ȋ{pi�NK�34��D6�> ;Q&k��%��^����G���~ҮF�\J��x�Y���?h��Tiw��'
�$�]�+��h�d����\)*Y�4�A����Kr-���ӎ<I�NRxP�w�z$��&�ݗ�/1�J��}b]�(W:�R��Z��[�_�	@�+q���*�� ����0J�I���w��h-G�׊��O9��T�It�g���P>���~��鿦7!����>�8������f��.���+	�-B�-w��nu��M�"��Gi�(�X�]*g�Gy�J�-�N+�?S�Q2D�}�J=�e��N�Ԙ,__��,p�xFji7Qd!/�ۀ�� ���!�W�I^��ܧ�����z闎H
g�Ѥs�5I���!�L���G}(�K�4m8�>y6��N��Ng@��G�b9�Y� ʧ��b�D
N;�Z����j�����T�����l�Q�8�ZG}&�/�'��e�2�{�2�e&WyO�i�ײF�>�O�y����J^ï�����j~��o�w��N~/���G�Q~���/�7���˾��ƘE���Q����$\/�n	wƴi<sn�pҷhs��
���Gc�1��6;%̍���ۯ���۔%���Ŷ�Ռď�В����߂φo/���G�	���~�,�k����<�� ��6*�0A�} ���&F�]lP�/��ȩv�{���$�-��K�7��[[.!h3<���x��)؟�&�[�$��{�)���i�7���W�+l���.�_�/�L����<~��e
��l�'X���	��b�N����]�n���=���ű�59�:����m���*���Y�s�s?�98d~珝?f�a��,�|��8ks��|��q���}����-��0�\�'�-}#cːk��wKZ�C��7"ߌ�yc�W�w#�E>�|��S��"?���?ic�4��Y���.��Yq��ǘ�ߔ��C���C��!�6ȵ2�<G ˳��%v����c���y��3���UP��������J���7��h�U�u^�׵�6��+ǎu��
���/ʧ[�|���s?�a��X��=�'116�m���w2�`�?��)��m��
	�Z�|�^� �<k|��uy֘+�5�g�5�Yc�|���԰�i�f?�s�'{]�9j�y:�X1s�ʯv����
������	d�|Y#�@��'���	d�|Y+�@��'�5�'�<ʑ��L�>���s�l�����ͬoju�¦֦���U4���"	��x=M�6@-Y�9%��YZ��g�D]����BB��3�vs�k�|�I�o]߲�|���R����k,e��O)�q�o�g��2�)��i2�s}��G�:��3
�B�ؘk�F���Xj\a��F���h6Z����Xo\k\o�l�f�al3�;���c�q�8hr�u~������+�)#�ЍD���n�9M���a5F�����D�L`�+��!��?BrR7�eF�Qc,3V�o����5�F�Fc��ŸӸ��a�2�5����ag���S�I���a��F������Bܭ�8u�`�^�^�]�3��6�}Œ���#|�������O����|��Xl\n\i�>#h�1�6�3n0n1�cl5�2�Ÿ���q��1�x��w矝�8�����O��pIF/g��o2���!>8ː3�Jd��)�\Y:j���Kzj5��Y��8j
�G�gFk�Ț�d�#���J?i��P�;V���TZl	J�Ɨ�/�c��Gl+��K��;]_{vd�u��M��
endstream
endobj
28 0 obj
<<
/Filter /FlateDecode
/Length 263
>>
stream
H�\��j�0�_E��P�:�F!JF!�}�l��JfXl�8���l+t0�-~��B�Y�=wF`�����(��]�Dp����a���Y8`Q�oK��3�����K���� ��+��Lp�j������h��i@���*f�e�NŸ�1j�2>7��3��6���	�^�	�>��@}��4�_�B�a��§l��$S��'���JDN�]�nD�,89�YQ͂��,)����>R�i��%���8�y<��޿�Y�T��
0 ���q
endstream
endobj
29 0 obj
<<
/Filter /FlateDecode
/Length 4567
>>
stream
H��W��$���+&^`�zW`,0ݞ	���0n`cm�����z�H��J]b;0.�Nm����!yH�~�bq/�����x%�}��ϋz����~��b��/�˿�rBZ��ܟ�y�q�����D��~����{�����vƪ���_� �����I���~j�o�>G���ǿ.o�����M	m_,�w:�Ň�o7���L���)��Q>~^�����@�O!��J��i�]�;�~3|�׏?5���h�"��	��S����u�!�B��!�愣�;+�5�Oy�Y�H�*f�Q�>�x� �����協M/�J�_��4<��h�=��"B�	������2�Q?�ӷB��zA彐�B���g��Q�`-�U��_�{��O��B<y��ۆ��8�g�����H >�m�O6�{W�ځ!�N��`�
��+�:ݡ6�%ٜo�\�t�GR�1�U��KK�N�
��JI��b����Z-�q�-�A�\����.%|���߬�W[�b!��F�I��O���k�����]�"�	��h�=LHR'�z}^['�Z����m��b4uq���P��8�o��GZ=�%�H�H˂�I��@$*�]0�O�'��&�H5��z���%�-k�+�jԢ�K;�0n�4(�H��=���U:�(t�T_\Ѻ�l����u+H�eѶ>N��T˰7�$ �����tºS�Z�[���.w~	(N�g���C�d��i9@I��M�KSxd�l'>�لM���G}]�4��b{b�2~�ݵ7����� �L���si;(ũ���8-뭕D����L�h�?��ە�BB-)h�R�\��!���v	���?�$6D�'a�H�E���9����ѭ:�c\��5�Vǈ?(�����F�ׁNx���vӿ��j��X��qO+�43����ƭ��栆�)�I�
�RjMoIy囖�&飥0U�t�Va �@!N� ��W�qȑ�͚7~B-)� ��#��;�_*V���o��a+aޏ�_�ܑ�v0�m����U��s*{$7�;X���C̩�J��-ٰt61���X^��1�Ѕ�?�4�4���)��TҝRz�U�B��RZ"d:��`J1�Ϩ��)�L!��=���sH����G7�[*�&#;�;�D�Fp�Ȱ���anrsH�c:����!��:,GӘ�D�-m��K�*��2ÎU�	m���E|:����NYW�O��g�w�E��%Y�n���[B��r���=y;��V��r.�;o�� r� I&��]��L��m
;��M�A��P�"�2�u�W8�Y�� <}@�t�
�͜�7Ҝ�6�y���5�V�0x�q������.������6��l���M�B���<����V�8L����To�D?���ҥ��{����X�D���#h���Ak���$n�q��[V�(�)���M�衛T�mV�H(>�v���-�9/���b����۲�-���t�o��=�<鴷%����\X�H6�L��>y�����m�N�&:��:UDj�vR�H���2G�T���VH����UR�K�L�t��9�a�:z���X��㜫�;�)��g�_
P�[�Ǯ{Mr��u�;?�(���(gD�ћ��.�<9ff�!����TQ��G�k����&�k���y��7C�Ҭ��Y�Ff��tj*r����]�dH~����(y��m ��G�<���lj	�"q�I���O aKz#I@ɘNm�%�`+%�I^
�λ[nU֦,Xe:ȸ�q�`�I�M~epG{��r+Q+anG+7�;�"Z*e\����U��[��ӑ ��V	b6җ�<�ڼ�v�����T �3)"OV�D�fZ^��B1;ٟ53�yh�&N�R���T�ٹ�*��y��}(�I�6��N�[���!mÕ�#a5�\&jxH�%�4v,?i��&�aZ�	m�=��O]NA*���Z�9Z�4�Z%-� �=��uX��`��8�#�(G�쨴k���r��=M�?&WZ��� �^@/�Z.B���;$�Fg��;�h�=��6�8��)^+ڣ��"�>˒�vk���x��I���g/����Y�;�3�����t��#�9sK��]q}�챻����sm�y�vؽ ���_��v���ھ3Yۙ)$Ԓ��4�%;�;�C��9��y5��(�}rIH�4�4	vP��'�'�V%������!$��ѵ�"14��n�����?D�qc�t
�t�"(��6��v���9'��893��ZR�����9D�A��rG��A'�X���9ZE��zw��L�W��_��v�Ж!Y��A!θ���D���*ŏ܃"4���F܃�BD�(h����ɹ�#�ȃ�A�z�{�Tϸ�|&��Q���v���6INy��m[�=��Μsd>��L ��r`�"�����"�V��eP���%��1�þ_����
�kV���c��tw��1��g\�	�j�j^#hS5�Eh�hwF#NKQ0���D5�$�W�صPǾK�|����nj#��!��~P;V��e؊ĕ$�l���3p�;��.�Ya�K;���K��� �������LѪ��#��G&x�"��+��o�D��юp��v'[���XH�4�s���+�ɥU���N��;N@�%4lq+�If�Ai�֗N)�%�`Ǽ@���T��;��z�Hx)G�R��`��%qD�%�J�)��2�`3ѷN��ǝ-<=n�9B�5��K��n�s�La�{���O!>br�@t������ ����m~g4��3SH�%�h
0��'p���:���<UR�H�u���OnW0�6�
ɰ�Ҥ3��Z��vtob�aK����D���/���`>�x�_ ���;�sXP��m �JmΈ�hFP��f��hdF0SȨm�f;�;�C�r��؁�ypFP�x��=ZI���<;�|&��؎_���tlK�kM�)��[�4�#�hR�s��e�.8�'�=��GF�=b��=u2odԢ4�&��8�'�3�0���'�	���~pz�8ejAЦ3�:�6&͙��h��)$Ԓ�^�\��C��!w5wqd�@t��sL��z�7�3ٷ�2�}� dkY݃B�r���WR������|���X�6�w;rG�Д;~2qG����9P����ku�Z�cߥt�|q��jB��C2����v�c�p�/��$�$���U����_y%�&g��/�;��2~�� �����x���=4�V#z9�^4�&:���v�;� w�d���)���㞳r%�A�4�aϘo	����V���$�4`�K��Β���^���Y��D�U]�S$������vI��*���k�n�x�O�`�����\��i/��A��%H�;���i�1Y3������zG�Ju��0nKug�|��ExB��⎗��?k\\GK�v�2��K<�xrt%�z>��z��;Oۻg�m�r$��-�*��o!�Y���0�rb%���6@�/�*H�?�]�3�oH�F7cU���9�7�{������3���Q}N%F�q݊��]�Q�/]���	�l�(2��C���,��
�R4ݮ7d��bT�l�OxN��>�������ӛF�G��y�/n���U�Jk%�g���u9�@���b>ΰe��
sh��.G�r]�р�0 
��zui=��>�1�pt<���������_�S<��%E9EE�R�BR4�(��Q�r$������,�}FQs +�`g^�K�+�M�ZG�de�T�q^�h����SG7^��v�{+���vQ`�`�!Y��oܒ�ij��*5�Q2�c�gH��ˑ���-���~���J�I}@�O8P>�gY",��}����2�ީ��"�&�ܩ�Y-_�V4?�R� Qd`�	X;����6h�tŸ����X�l젊�j���T�6wPU����(x�j<� ����A�V^�%	9E�ɸ|�E"����C:^�$4� �؂3�{������ф���D�u4 +���xx�Bԥ��B�O��v�>�n|!Z�K���9�8E���Q`_3�q�T ��H0cU����`�>��g���
r`��TYi4��� ��z0}bC�u����m�`��
`�/�$��' c� v9 ���b>M f��
sh��.G�r`�р�0`
���ui= �Abc���� ;�� �U ��"���w�� ���r$g�N;��V��t�������o�z���4�q��7��<��N>�-�������g;���jx�����e�Ȃ&`܋�ed��*��,J�g�q����t��Ѧ��C=m��ep�UU6qnbpG}�������������I%��G��������޹:�*�)$穻����U��E��/>�VƐ�|u����j�.����ȋ�>����+g5?��9��7�g<-[�F����i�U��c%��/#�9��D����.�_	9K� �ܹ�
endstream
endobj
3 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 4 0 R
/C2_0 13 0 R
/C2_1 21 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents 29 0 R
/Parent 2 0 R
>>
endobj
30 0 obj
<<
/Title (1ec8b7e24be6c30b4bdaf70cc209ff749bbf40476b630bec24ca6359b02604cc.pdf)
/Count 2
/First 31 0 R
/Last 31 0 R
/Parent 36 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [3 0 R]
/Count 1
>>
endobj
36 0 obj
<<
/Count 3
/First 30 0 R
/Last 30 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/Outlines 36 0 R
>>
endobj
35 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227170051Z)
>>
endobj
8 0 obj
<<
/Type /ObjStm
/N 21
/First 157
/Filter /FlateDecode
/Length 2675
>>
stream
x��Zko�F��_1��=C��4��@���i���j�uؖa+�����{I��I�N�.� �������̸k��M�$S|,&�H�8��V�p;4�qٔh�q�G٠θ`���xoj�(�;o|DY����dQ��x��A��46��(����j�d�J�}��l�ϛ������<;:[^mV���g�����W���l��w��\__,/Q��ً����g�nj3��p��x�1�b�?�����ru�����f�WK�z���__,�oM���ڼ|���99�����A�l�T�^\�.0�WW����p�~�>X],�qN����˥�|��_?��N�����bq�u�77���������rq�7?�H��؎6����ë�%&:?�,/��g�_��:�s27���m���e�����������z������6E�����1�v����/�ndx�58��q��̉5'�P�|yP�!
�PY��,�`K"��
<����y�O������)��8ܫ&g�;��Q���ٿCa%��������2�*�Mvm`�.��=�:[�%a�Z&����&0<��c�ɳL��*"ǁw=J�9G��o��%�'������B.&X�M�`\�&C닰��-���s�Rt	�w�q������'b�����q�^����96��>�/ ^ b�MA;6��A�'��/�@8�r��bT*&-�ᇁ�)�,Q���Gv:��Vr���~'�2�n�{���w�_�r�X/$ܜ�i���,C�0B��,-aH�Q�l I����$!A���$I��"пC/c��|�"g_Tǜ;��{ْ���&`�^N�P¦$��6g�P��9@�Bpdж<p�B� g�?�ZT�+�RL����W|p6�8`4	o��H��u�G �y�J��(`z����
b%ٲܧ7���U��w/�m�XR��,������p��DE{�I��UFٵ'uX���J`ܭ�T�s���t({�^ $�>�)�Ԙ�xUz �A>���ރQ���o�k�1� �����F\6'V�c�-D����7J�Z�SW�Kl쥤i����TГx���f���p��� ���*�u0	9˞�������.��[��wiC������5,NyLga��V��؇�ɩ� G+e�+ȕ��*LdX1|�s���HU�n�9$6"�1�u��y���Ϊ��$����Zi��5�^�xY\'��꣎K<������H��d �S���!zyLw9M�pՈ���%y����ls�-�Vf.��6̵����ח?��'����.S�E�5�6��~�ͨ�(�.��c'�����.j[J���,l�����6 �m76^���ħ�~׭�� u�c�1m/ʽ~�����w�w �s/��{��<Z0�
�!ۋ�]̝D�ʌ�}H�@BZf��K7Y� ����vJ���mW"���`��B#L���.��f�Z(-nW<!��p��d�޲�6�ށﲮ�/Ӊ.>��!��7�v<؄�o���ǆ�����r������H��G����*~
�ˮH��d�2VA9�=w��J<�MS�M�����"!�0I�B�&i���:&�A�Br5�m���}"C�}Gpqȥ]�Ӑ,� iR�w*If�I����åA�Oy�VI�Cm
2�(+��C�T5���=�Ç��>G�����w
c��������p�����7����q=��)�u!|��z=Tn �<5�&���-��t��):���6�i_g�}��s�e�t=Q�>��n�0���`_XS0MMI�K����p�QWߙ�4 SE:����&bZ+�S]��V�b)}s-�K/��$
�Ю�eG�	�&7L��2�]>E���n�E<��`�r��'���+��	[��b�8oW�$g�6�@��{�L Y%#&��y9�.����gDG�N��d�M�d@��D�sЭ��E�o�L�(�$�uF�xB�����f���@SNJ��}tY�0�n{�l�<��Ʋ�}x(#�2��Y��q���c�7f�������ݧn�)�p�{M�:��c�U���-���I����|��y.�}����s�I��+#H9��޷���;j�7\eS1�����$��tp
vx���/��N��T�lq�a�[����W��g<��w'�o{�_ݹ���*.� ��N�0��qfw�yr�@y�][
���3�$�rG�\Ur�D�K$�W�sU*�DjxQ�6����ڊ�K��K��K��K$n4��<�*/�^��٬}�������&*�,c�������jm�������t*1�Q��[��ՉJ��H��D��GgI�X���w�2�:�B����%�\"q�K%�*q9��*��@$&h{�[N*�%s+�/�2/����R�%R�K��ez�^��Lof�{��s�d���a�Ι��J��y�K�a��q<��~s��������;J����sL�4�cz���1��w��<����3=L��y`��uNe�������xq�t���vcƴ�p0��H&)�O)��R�(o�?���CJ�4I)?A)��J��(u��ݿ������54aND�x�ڼ��ʧO�s����>VL�ٻ×%�g��j8�v�]u?^���Ԇu�^��n�?AR�ݢ��k�vM��i��
endstream
endobj
37 0 obj
<<
/Size 38
/Root 1 0 R
/Info 35 0 R
/ID [<5217C64AF857029729064CF134102380> <95A05ACB0FB41DF3E42726DB5476C82A>]
/Type /XRef
/W [1 2 2]
/Filter /FlateDecode
/Index [0 38]
/Length 124
>>
stream
x�%λ�``;�<��.̂�D�h�,)C	;��騳 ���u�'�,� N+��j| D����8_� �XDo��
��HY/2��v�؊R�D��ËZ4|���ӌ��؋�8p��i,'�-;
endstream
endobj
startxref
49463
%%EOF
