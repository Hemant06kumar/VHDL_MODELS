%PDF-1.7
%����
10 0 obj
<<
/Filter /FlateDecode
/Length 22
>>
stream
H�:��"������� ` 
endstream
endobj
11 0 obj
<<
/Filter /FlateDecode
/Length 2248
/Subtype /CIDFontType0C
>>
stream
H�|TyTS�~1&7V��&��V*��}���Ȣ�� @X�0	�
�B$+�"�P��[��R:�Stt�LG�::����}���/L��9=������~����w�l���`|�us̎���R���m��c%�y�b�7���S�F5�A͜J	|x�<����q���g��K�@���8-�'c�16���3|�6��ɒ�T�L)U���Eriz�R�x���^\<�K&1l�O��%�����d�D��DqE
�$G!�����\R.VJR�6dg�&K+Dr�B"��N�܎H�I���\$���RZ/����rq�$G,����Ѵ���H*ѵD;dR/�Sғ
�X�BW!'WI!�dJ�T�X�).�(W"Z!J������`�F�a<����~�-a+�O�MX$��`q�l'��I�����z��b���c>�fʜ)}�y̛S���� k5�4۟��~
�g�W��2h�ʤ�=�nԊ	�Cv��Y�s����^��28ɐ�Q^�ͤ�+�{n0��	�<T�.�g�B6���:�P�5��p�P��>NPM >o{aT)G	.W�.T�u	���u�P� x�0x�
��ݏ��^��7L�� 8�[��pHX"��0Z �]`�Mo%����;��}��g�*6�T���͸�2!�
�e)���6EW��q�[і%<�Y��r��t)ڳ����Kȅ��^��iğP�?0�����C�]������ڥZz�2 }l�B�p��3�C�ʸ���V�B'��hJ��t��&��8-���C*�E᣽g�(l)�O7f�x �5v��ao��!;���c��ϧ��2^IJ��P�`�^�ߝq��PXT�m `�w�M^'��2���z1!,`���:%x�wi��uy5y��N�L�5�X;�e�=$�Rc7,&<s�*��s<���A���W�n����A��������W�Q��Xl)�?�x�����]��L�[�_����*�,��d�(���Q@1J���T�ݯ�ЈJc4��w���Vq��w��9��x�UņJ�)V3��,3��Ypt�^�J�!	��y���`@���/�����d�kQYS9�l�8�X��}��Q�¥X�ۭn��Ւ�����д��o'	�����wF[._7=�� ���:or	,�m���.���\���X���k�|p�#ڄM6eC�����?{�=��Iwr�։��^?�H0�����ܓ�(��?*�<⬪�m��$�����\dO������P`B�"��?�I�Kb��IE`�]W�8�u�����#�/~ܞ|"SSM[���F��1��~I�K�3�P��)�;���^��/��J3k,�	�H+�r$A�Q�q��A��h6�{�J����1���n|T벶�	�{Y� '�Z��k5s�^r�W�H?�Ώ�8�ù��]:�8�!�JTc0���a�q�=O���;�4]r8���ڛ0�R���5�&N��bo&��rEܤdA�>��Mb�������������ĄJa�V[$�������p��%>%��ڂ�o���܍��T7����:��J�*�rr
�	�y�yNe�X���_��d��n�v�IM�d�Y�ݪ\�ftNl,`<u3ay�W���!��@��>���5#:�a3�����#�&]�oo3��a�7L����s���q��^���6WD�]^I����km��
�i\e����ӿ��ď�SU�++���]��]�{ß�+.|�Tr�-O�1:�����
�^��a���� $��W�Qs���ڢ� P
��h��]�CN�Ϊ�{�;a���u��?^�=R/ć����Z�Du]s3A[&M<�;G�EKT��]�^��;Y�be��/�l�Jk�jm���b�Y�����$�+3����5=)#���Ս�j$=���kk*�=���MT�YŒT�mW	���v�&���?^f���dJ%G���8�	!pӘq�tJ�K,O���f�����6�<�j�7v
�m�mMm������/��p����í�/K@���F<�΀�R8I��9o������y3����6�s�{���,��� o����Jr����ykyjwlwnP�y�������\r���Z��n^pcoh�cY��M�q�O�W�������������	�p��`�q 
�&�	[|��I����%���������F�_	��
��w�c ��D
endstream
endobj
12 0 obj
<<
/Filter /FlateDecode
/Length 303
>>
stream
H�\��j�0����\/J��B�k7��,�����8�E�~�T:����_�Iɱ95�H���Z��=N��+�3^�Yڨp#z��9���v���GQU�|Dq
~���ϸɛ�荽��ױ]A�^���m��4���K�^�!��u��n¼�9��Cȉ36�F�����^PTi<5T������g��ν��<�g1<M�^(ˉ6�d*��D�Qq"�l��d�3�
ֶ��=Ӊ�H$�K�^�)gb/%{�\�䚒�+w�򭷥��#�OV]��C�E�4�9��]��A�Z��` ��
endstream
endobj
17 0 obj
<<
/Filter /FlateDecode
/Length 23553
/Length1 50984
/Type /Stream
>>
stream
x��	\U��?����9p@Pp��#�<% �("*�� S����sZ��yӼ�f^_�z�Fjj�e��յ�����vͺ���k�}���}��������<���^{�g=�z���B	!~��LJ�S�����fGo�	�I�߫(#d�z��66#�y�!+b	xkDƸ�)��?J��@p	Oc�ԭ:H݃��s��ˆ'~�P��̮t^�� w��	a��e3�'��?%����}3���@�?�{�̢y��~�BH�@BB��e�Z\�i��+@���a<��}���ʹɎܸm;��4'���������}nq��2�]��0~8K�����J"!3;�vhYiE�k	���>gYy^٠�N ��<!�vRVlj���F|5�g������wO���}�yU=U�Y��x(~0�R�w��.��������(�ǫ�&\�3� [u֕8��t=Q��[݂�`���'��<5nUS�F:��!��2�*&��'�X�t�4ݟn��/����S��ER`^ea
M���H�t/�Bv�,����k$�,#��f��uh�&K�"z�n Yn�v$�Wc�"Ư$�H1���x�V��
3W�(���a�6�6ɧ��Hp�X_!���)Y�ä�� �S�s�����e�{����7�ǐ��X���j�&	G�kt0z�9�c�P��x�D?��Y�{54���Z� �Ι`�<�a�7���GA{#t3�pЄ��7dA
�L( g�����FoӲx�(g�P�[�'I��`��r�� ��S8ɾ�X\� Ѧ���S�ueCI��:�`u��j)��ݸ��{�"~�%�۠=w9��a=�`�!d*8����
i9+�0��Cړ8��i��OI�F��',m ��NR3��n�ǃt!��V�������=��I��q:��b\�_�K�x'��7h�@φ�k$$���C��+�w�9bj툩����@JԽ�[��~���-BN���T+��� �0�0��+eE��/cV�`��� ���\c��|@0y0�����|p����y��л>� 0t� �j"ًz3 ���; �Q�-`64�2���$>(����xR����E���^�n�����ؓ����?���+�!t�랡q�����42��m��)`*���:ѡ��y�C ����F1J��]�#�ҟ��hO�~���.]K����#
�!f�j�i������L�Ú������ަ3�kڷ�!9o-�O���#o	��\�?Yd-�(b��qr�j�'B�S��|}%l�K]���c�a$�^suԿuut�Y/s�E�I��>�3�a�E����J����`EU���N��Oano���wV�~��5�%	hU���M�~h;F����g���R�܄Q�z	�>��)V[M���'d:y�7��a<�	8��ՠm��j�Ӻ��~�;���-	E��T 9�-��H�+�R��͝8S
H<�K�}9��wF��옅�"���d��P�*�:%���s0�A�K0�ŸT�G�0�?��tP�I6`�Sr���c�8�%�>XIHT���dy X�?��J�d�,~Xo�Ι�k%5衯5�1�~�/�o[��z���FAO�l?'ǈ�9d1h�z:lc1遻���o��i��G�E�����0]>�7�9���F`g�G���<��(�Ë$:؅�m��q=JG�������l;)�(��}�|�{`)/�7`���?q���]�H����0	��=�!�+� %�e�����A��$�Q���k�y@'��倦l�#�j]��+N�@�A�G	M ;xS�7A�B#���`'9K�a�'�jb0V͒k���u���Vs~���y��$٤:}Z�EFKO��8�$�Ka3���8���^E~W�*�0 �n.It�`���4�캁�v��q"��קͫ(�e[��q:��w�刧1�i�|���fk5�ݏ�����'a�A����
X�0�:��HD�A��T��DڎD���RF��U�%B�?��^���4��睌�Y(��3�N&.�ё�iY@�����,��A�7�u����0��c҇0+\��I\��\:�\�NDz�9�{��K"�pwT�.�k���Ƹ#*w�tV�={�ܱFy�y,�7��ќ᳎�bDS���ע�;ETa)e$���[DqA�8K������;�p������������#�3JR@D��E�v.���:k��Z�ZT��~�n������S�U�^��s���!>��v��p�v�sw��s����&��J��&ާ�U�R�@���z`K:1'_�yQ���O�K�g�</���{�S/�_��/x���n�ݵ+�~ǂw��F��ZD��oA��MG���r�S���#�@f28WA�d��0~��݈-v��"�q|wGC�Ml�"��Q��s�X��45�죭�b��Dw�ȿ��(fM©��7d�6��1/�����%| �C�����y"<� x�^9 �<W�1��+/��&��bԆ�p�Q8�#��	NIذ�����L�(9>����q/����96��=�}C�1!0��L��vߙ� NO����A�8o�6F�:��rF��V|S��<eBÓ&�DO��4�xy���%V9ZQ�1Q���6Yxجo˼`��7��=`	�%ƙ�3Y�.����ȉ�үQgA��'���f�Q���1c�	~��Y-�~	K��T��_@�	-g��s�5DY��\?!��dґ��5��i2�z�b����(�;�`W���)��QD�_�ѐweQ"�5�X��u��7y���� �]Ds��~B�Ы�qS.js5��_���6ٗ��g��V��m4(!�ݢAf;���b'�̎��<Q(,N#��ղ@z����W(jzV<7�������]��UK��:��u�{��/�������H�f�m`���u�*I��I�v� ��H�e_����T��&�D��2f4{>��_�O��g#�~�P�t(<h��A�,<J�E~��#�Y;��w8푽�?�"�>];"+0�"������g&��Èv�4�1���q@ v�~d)����!�
��@� <�_0����z̛j6�/�s6�+o`�Af�k/I�q6�"���!��;
�3Yw'd	���Dd	�"��4�H���+tAV�YS+�>0~:%��?@�9t���J�A�=��:�F�f�X�Ln)"�X�>g�S�U��:x�c���lÑ�G	C�	�&`L'<����hE���X'�րp<q�7�n�m�:�+���I֎����c�.��-H�/	O<7��OK�'�w o���9@2�R)KO����dN4]���H?:�ȣ�B�qv����������r:K
�'��U��J����ȵM�|��X��ji���f�<qhD��;X�:�v<�ϒ�B�xgN�����6dYn�L6�7!�f��ǔ�����
�0ڿ�a�_��\	턉�Z����:���*3�߸"ǝ.
����~�����qLO�zP��Qx��*�;�h��("�'�O�*d4�b�����Sh��|���ίp��� )r_���WDl�ͮ��Ʀ��tt}+�V�3�:����d��7��
~/n~\�\�$����4�'���;�>5�}Rr��o>D$�!2�y�3�o'�Y�v�P���9�0�Z�j�u�j�<	�tl|"߄�>�X>a
(}E�SQ�'\2'��I=�^*��ٯ�bgx���3�x(|R2�kV�)���&�h���˅�b\`�ø�K7�e�"x��G].ח�N:>��'t��c���}3�)��4E�j���-��|���_�8�(�P��!5F��x7L��Qb���O����c�F�d�w�Y�Q�QD<��R�Rf�*G�m⚋2e2t��(8=�ϐ�� ��X�-��_H�ʏ[�#��c��<�NDC�>ā���?N��8/a=mqζ���}9�9�`��!Ϯ�gwbHK�)ڔ��M?�Ed{�)�'^J"1�D��8�FKI���fH�Y�D)�)����/<��o��h�T�#�p:������f9�N�����8��^�5.WZ��N�x@m��[(�a�����{F�N�r��6�	&���	���BSܡ��	�X�����8s
�����r���[Ln�O�kOpXsԋ�B���v+Y���8��m��}�V�޲�u��#Ըp���S;̌SO��6��C��"���"ۚ�ʶ"���a���NԹ�����N�?��v����B��5�:��r뇉�5��b凛��&�b����?��R�q���K�7t�]��Ͽ��kAb��kk\c]��G�o���l��r��:��W�Կ���v��:�z?�R�_��~~��?��?���:��� �#���l�� @���?X�~��_���/��� ~I��cS���;6~Q�t��*_�������M�����X�����u~n!?���t����l�RO����O���� �����{��zL�/�O}�y�r�H�z�>~4V9����M�f]�����r�6�3p���?�������^����z��:ߧ�?��:n���\��͟��>ە�������������:ߩ�gt�c{��#�oڡn�O;��l|�Ο�"O�|�߲9Rݢ�͑��Wo⛞<�n�����'��'+ׇ���c�:B����#|}8_a��㏁����ZO�kr�jmu8_��W�|�Η���e��:_����R�?��>����|�\�衅�"�?��/��|�7���9:���J�Z�ëj(���T�y�	�W�*�:@�e:/-�PK7��jI/�ʋt~����^p��<��u���\���Vst>�8��<[��u>M�S'y�S��}�|�Y>7���$O����t>^�����bx��3t���{�4����:C{�ct�r����G%������~jr �����܍��I�K:�y:�����p?>����z(�q>j�/��awq��j����'p;̮�z���w���0;VCccs�{t>$�͇�|pW>H�!���|@���Ѽ�����W���h�'���g4�Ko��``��{�q��<�-�B+*�Gz�V#���Ԟ��g�F8|ՈV<B��I��=\����=�wc��n:��.:����[ǫቼ��y�����gO5d!w��G�`���:oٶ�y;h�]o�� ��0�I�z���y��C����Ƶ��~��s_p��X�����|���1d��eS���ې�d�e�^���݃ۅm�W<un'6�{��V��\jM�?�`�����Se�8�''Nkh���;?����?�A�/�^�8��D�,g���A�����q5���F{7�C��|Om�5�K�Y �TBлف�����T��]�-��7:�c.}���O�me�*\|�
�~�g!�(&��~`\�5K�"�+K�7�o�!�_�@v�R�eKA����.7�fv��{΀ǯ\�^F����eCY��݂u8�ҥȆ*��\'���Y`}2�lS/���<p����B:h5��%\��Gi/�JޥⓄL>�?�?�˔0e�F�1§#�[����u�0�N˧����e:�K����C��j�	y����j*xΗ��$�uF�9ț�6��8��H%�Ó�x������u)��K�u�d/����o~)ڛ!�c�t5��i�������z�,�/�nbYH*T���"�/�7)�.���񨌣� �CԪ.ENu�Rm/�T{�6��o�ox�oH�B�*x����,�?}_���I�{9d+qu��+��J�)�(>�n�����a�������'Qe���8�^�d��يC�p�Ǝ�Ě��տ�U��"c}�m�)o/�~	�yc^L�����\WM5���&�3��ǯ?�Z�t��7Vk~W��_�U��uz�O��Z���]�x-��zZI���	�u�1�x{���g��~~}�0:E���_�>����!�_�W��J_�n�?g��(�F�����d��ځhB���xX+z��������.2xͥ��b���=Dv0����N4	��̣�G�t�^�B�����ɰ�!�(��7�^������^��W�K��&��`�"�nJ�7���]?�^�g1F.s}��`y"���ض�?<����Ձ���t
n���v�>�!;�'�q\��7q�t=:��("�@D�(%J�Ң,Q�(�([��02�c��0e�:Lff�1�6�s,Kǲ������4:�M�M��N���l;߮lW�k�-ۭ�=�۶{>O��ϳ�����������{<o{��89N�����r\=����8n;��kĘK�i�4u�6�2�:�C,�k�:�G�}���i௅�vn�|~�c�|����d�rL�ic�l���k[����~���n�d�������¶��s���M���4z�>W_�?�ϥ+�Ct���f�]O�$��F:���j�U�+,����sh�J<]'sSlbl`�oxo_a/�t�����N�՝ݫT�Ԍ�}y��5���A��ɽ��H�pUS���6��5M�w�>�U�I!Ռ8l�ڂۄ:x��:�uℯ�@s��磑�Y귾m�K�����X�/R�{h�>��B5K�{h�2�xSZ���U��}s�6,�|�l�k�Rω�.�ݻ���g~�؅��?�+����OTƉ_�&+a��AoW2��������U�u\��ݾ:l��%�n�[����C;�{t�zA�Z묅y
�u�q}`4��
�إo0��Z{оF��ܺa���f�73���ܼu��m�?:�X�����Pu%���'��{�N���ٴ��-��W,�������쒾S��J)���q�c;R/�E8��'��R�R��m$تh>�Nގ��KC�������@C��9���P�{��N6�/�T�F������/W;����Y�{�����[�������P�ҡm��w��1�j/VMVxm�����M0��G�`����~�j�K?
ZA��B*$��4�����f��"�����I�r8��?y�ޭ�߽����7����͘^v�8i��L ���,��m��?(8�S�[orl	&��B-Z{ڪc�p7uWko���:}�πH*�� P8�0'�"	�iMC� �����a��9�j�ޒ����^�=���6�/ٸqɣ+V�/���-�~��|�ߢU�q:���X_tx׮������Y}
�����Aj8㌇+��B�\�T�������I��Z�Feb(d��CV�}�߼ˬ�}���o/Q{�7kK!�T�{�Hh'�]�����~�]���w��)��#8�](�	���J�	i��]��l�� <���astBO+� (�,�����__���.~���M�u��Uݵ}��y�/Z0o1;S�jՖ�5+7g�����ŋ�rv��W�<���1�����_�İ�E�)I�ԉ�m����px��?�ժ�o
��J�c�G��s�P��Zh�}���Zv�~��??_o�w���~B㡝Y����m�����'T�^�X�{�F�ɭ���P7�A��S�����*�T_�Wt�<c�.2�i��v�}�NM��p�R8��Ɓ�k�uuJ��>P��!��P�	�meE< ��}6����A�!� ���j5�.���'�%�������Ze�2��*������B�tF#�����h@�Re^�~���JE?��z���Mw
�d���<���Ѯ���bU���阆�P�}��ϟ2�>�W�6{a��m6�96��#pY�bA��UU��6+
�q	G��m�}�jz �O��Z4���C��y:>��:j�v|V�o,ƿ&-+��A���ض6�#�\�ԓ)ܮxX4�t%��G�<D9!<�\F\��蹋%�?]T����v�L_ ��n�� ��_�^)�T�<��V�j�;�zulee*�n�ƴ��A���C��͓F��Zy��^}�M�ݍ�&[��|w`��{���K�l�G���i������I�\���>������-| w��^���w���A�S����Hdl۠?�����ן�������b줗�V���.���ñc����mL�)�~��^cvN�?�O�a���cF����3Y�%��֍n�e��n����_����/��6�2K7e�56@��XA�}4��a�1�^�`G���! l�pg?_G�0�V��nԗ�@\��s��t<MЏ�{����#����F������E�E�'/çt�m����H��GU=zYp���K��>ݠ�;��]���/g���3*io��f|���d����ĭ�C"�c3|4Ev���Oay�O�!0��[�ߌ��TҠ�dHlHP[Қ��n�L_�킂�_��o���i��T�~�:b.��_לoX�%��7f�W��4�v��/�޽�Μ9���n�[�C�i�P`�~o�I�߆���;���wKρgM���&��T��������.�:��!�i`�/�s|��Xw��_�?/ڻWYb��}��ȉ�R�4��"}4�t�QW�^d����b]�zYF���Ǽy�g'�b#�8b-�3eԃ1o�0N����	�ߡ�4M��i$��04Ç�ƜF�<|��;�:�c���N���ц�6�@�δ�l��я���<�}, G��*a\=n߰��y�#��-����Z�O�{�]��n�{�
:��Ρb[yT���M>[I�����7P�>⢩;��֪I��\�u���[�.����[?�!	�F�i[�+�E�F���d}��y�
��.��=�N�o@ȯ��Y��d�M�
W���k
	�J@�������C�6�K�{s[P�����l��`�����@Y	��\�o��Ƹ�[$CX�i�#i�χ�����RK�����1r^y��E�g�/|��c���+����:���W��?yg�6���Ï.Yi��Q�e�H�P/;���l�`[xǎ��6���
�����վ�O�Y�:|��6ώ�,�s��޽�-C�������*��tD�n��L��d�d砕���f!
��0*N��D��yD1V'�X�攗���]��wN�?�^���͂-{�/�p�z}:������C�=�S��?_��g���V.(���:���u�Q��N��B��zk�/4Ho]d�װ!�(�B�������e�x�B6@~Ce�-���#
����+�}�}{�`�`���B����n#�ɜ�)��5�nx���7~��������*�;<q�7�ً�<d��)E�V]�__6xР���1h�?Ǥ�y5v�G������).V$����p��S��g�ē"������8����բ�VkQd�-��j�Նmߦ�eZ�m� Z�C���p�T�3P�B��njg�,Ϲl�:��S�����X�Y[kb��pϾl�h���c�!Co�a�G���U�_�8��_�'��+�&\Û�w}|�5��~!o#d�2x\�/���F�`�Z�"�V�רE�h���|��fI�A��)�D>!\19�����u�������?��ݪ<.?��;(u�v��Ϥ!�:o�]�L���QzqZ����,LY �VR����i���C��5~!���;��t�oK�T��m�=��h�tG؉�c�?�:}�f�M3'�������1����;��ϝ�w���#hG[��̍%���8֤�!AL��Mgd��.ٱ���~~�������i����������$k�������eye��R�dw�Wv9���y���t钞���������$:�m�݃���X���X�����߈@���M� �bb��-�c���ʝ��^*sO��s�����]���e+꿌x*�������%���E�w��˗>���g��N��~fB�Z����S�'�"Q�m�N8����p��c"��-����iw\��o����[�J��ߥ�u��4�*�nMM�p�>�o�渁=z��0�{�+q�>�����rY :�@�Ð�J�ۮ��_c��}�>��(Dc#|�<G
��7��Ȉ��S�5m�_�I55�[r߸���y[u�˖�^�l�
~��g�ڌ	t0@0����ޕ�.]�����,�% �$�vFEm�=�j�Qm�}%hM�c^[:p����Z#���&m���7DuU���uN��M��%Z3S��<�?�Dq�������ޏ5��+��s������"�7���v�rf�s�	�aow��Z�>���ڭ�4��<孝��V$9�����ȯ�bɍr5F$1~BrX�5�y���+].挡K�E5�e��?i�[��.�_\�Z�߰��H��ܳ#c�ك�u��~�[��X�z�ǎ�9��d�.AD�����BFbÞ6��z���Y�E�9��}��g���P�D�m��擖/Y�غ���\�[��;�?�"bs��o�9]�)��|����~�/W������EF�<`]8u
D-�J����q>��������74���?��O#�������^�[qH�<��Obe:.����Y,Y]S�kO��c��G�CՏ��������9���z	Xσx!�
�"�Ӷ��I�Rx�'��2�f�®��1^���zC ��=��>-�+����cM�2�.j�:φ_|��:6�#V�h�p�!�~H��4��yF�y���<)[f����}��E�'��?����~J7=�жK'�?�o�x������v	���P,�C;�`_���ڝrX���u���;�'�}����a����3G�͜��i�:1`b�6�w�C�\�)_@�
Ď�V��h-�m����E{k=�Ͱ�aA��k7���Â���bu��زغ�c�m����ڬ\���v�گ�.8��'�d� �DY�Z�ٮ��Q�K��MJ�g���>�3,%�_�xQ��~[�mł��/bKn���2}��aI�Y����w���w���a;��=�tD��4R�9�kk���8=�|�_�=��5��M��5�Ȁ�Y�~�����^���7�n��^y��^~��6�����ҞTD��b�c�x%�
��;�}�o>潅��';�/���ɩ�������4ϫf�؜�^��o_�����Xn�a��֟�l�2&�����:7��`c��W� ���ɗ��$,����j�c'-H͈��q��Aĥ�´�c��A�N�N�hM{;�}cI,��M#i4͑��w5��FݴQ������<�4av?>/�����U�8gQh'Ï\�n4�ӅT��ʜ���2�A��!8Pfd5=���8��WY~iC#m�N�N�h���]7�,mp�?�Sׯ�k���D�E��5M���=,s쎌���8j���w2͚y4s��?X�?q��I���/DFޛ1zT�w�mw	;ַo��Ž�w���y>D����O��{�z�V~��ғ�C6���!8����8�7���s���Y�����|�S�:������+��i����ذ�6}�ǌS�)S[�-6z�.��(l8�׌wfV�N+�B�Χj�/{x�K/�z�}{����Vc�~޹';�sC���X�N4����6F~І3�PYk񌓓H"�%�$Z�{P��D�]d�-<+�*���s��4,�8M�I���o��3���w��в�x��bG�m4����E\T�2��0F=�`���������G+�|�E��t2�Œ�Z�6Vw�L`���	�E�����%�Zf�y��E��)}l���6+��`a2I[�T���\�k��.���<�F�(�뿮������H��O�4�^ _������^m�����<����̷��s��qq�uxy{������w��"�k,�|�O��u�x������J$	�gr�*6{�МW��˷���[^�1����V� {�Wg��>|�}��&z�D^�Y2Tー��S�%�#rB#WM�X|���S4��8E���?JM�:���Z����X �z��X?Df`� ����چO[���MN~��/χ0�9b�h>5���Gk��}Ȧ�Q�i���îy(^0_����j������Fv+�B#z��U�.�3&�u1cE)�߸��[����f�9c؆=���9ċ~����1���b���6�@�c�?�m;d�V�'�T	�`cyxZpt�$�z%��dI���)d4Ʈ&5J��^��Z��Y�. 1k�PҹF6�t������Z���3fg��4��4��_���VN(ߨ5Ƅ��u��V�m�N[Z�%L�����/<�Q�{��i����g�g��a�[�I�'�J��k���Z�~���o�D�������ul��8q��]�w�.܅�p��]�w�.܅�p��]�w��>�u�fޅ���O �����hq�%#J�3ڌ(���/5�+M�*��
��o��l�����l{��i��屁�c��I������1[�٦��f��z7ۼI�Ҥ��@��f[#�=s̶��z.2۞d��3f۫Ug����&��/-�W^8����5��3&:��s�<g|aeEey^vq�3�$'�WT�L�*��yy��r#m	y���W9s
�Kf�U8���%β�E�9����������
�Ғ�������W��8c"{�7����9:��Ub���ʲAQQ��]YQZU���_Z>3/�$�2jN���Q�%�ys#�
ʢR
s�J*��lA�ਁg׊�<猼��9�"���6[�dМ�407H���7l���l�-V.�����ܼ�������-��liy�ŅR�]�W���f�g�T��F8���<��aH/�YY��.��,�*0�tF%.,��Ur@�YY�g*";'����ŀ�`/2$��*E��r���9��X̩*�+�̮��A�]F9��Q�_92�&))�++/ͭ�ɓhr�Xጪ�<IC�	�RNQU��dNaeAiU%�).4��QmU�v"��y�k�ߊ��&kD�5�J˝y�F�T��K‶L���\hNAi�/'5�W��`�<91��YQᬨ�1+/�R�2.�I
�rJKr�l�L<ʞQ:;Or`X�$��JJ+��
�Wh����gΊ�l05#ϔȀ�g7㳴vQ�,.-ϻ#���yey��X(� �����yqina~�0��J�@���+97D'�Wv9�*�.���U�,�d�,�WVP!&	���
1�MOE˕��5�]�A$�<7-�AbI�<ga3SK�y���XѨ��qo�<�]�������
gh�^k�8C���b�vL�Z���*�A01���������5��2l��Ey��?0�PLAv�� ��J���5Zx��
.Ҡ+��_	58�-�V���-U'��,��=�,;���`{��������l)8-��W�/���L������9!.=љ��LK;>9!1�������̑c�e:1"=.5s�sl�3.u�strjB�31+-=1#�96ݙ<&-%9}ɩ�S�%$��p�c^��LgJ��L �+����3�1���G�6.>9%9sb�3)93U�L�8gZ\zf��q)q�δq�ic3�#hS�S�ұJ�D0D�ǦMLO123�2���L�KH�>:BP8,�;�HP	���br�ȸ�g|rfFfzb�1VHgD��1BF�R�2�Ǧ:��J\|J�AX��<&7&nDbF�"b��N�8Ą����q)Ό���ɢ9&�'ϔ#!{H"E�;|ljF��Ёq�%����r	0��%e��T�+�d�M�l eBrFb�3.=9C���>�
}b��q�)��j�+t$�~i%f�&$ƥ a� �ca]�ss��*�m���p�ҕ�3BZ��`�#J�q�>ل=cgɓ��p��K����֍��p�����+�+��(�dNa���8�K�s�"��aV�(���"L�h ���r�e兘2����ę]������Q\nU-9����<��'U�켢y�[.�3IIa	��b�u)���AnZ�)��q�j�N�`���#夐�$��8IW�C��C��њ�N�1��+1:�d�b��dR���k�� N�ހ�B��ᚇ9�Q�b��$�5Ɠ*����l`�)G:����R��cf o!�91��f�g-�dH,��*A�G)%��X��J%�Pћ�o6�=�=�9�|�kpTir/8�}��<�5����H�+ŵ\~Ր�[.���<̉"s@��(Q�1w.��g�R$�y��<��dm�l�:��Nĳ
������ �R��Mj���#��z�ieC��h5���6f�v�
b��v��<�Rt���R��R����v�h��I|�[����<���r�i��O�|�װ��a��"$]���9����
�k�*MJ�0x�1%��Y)�h�#��j	)3��1���E�lZh+����J�e˽��_�U!�\�m�?�s`��K�|�O>ZE�wm��q�������e"z�P�b�*Ig#5���Jik3�R>u���+D�{)�UI,�L�H(��ҔL��kʑy3�4���2�h��.��t�q�V`vį���g��RN����BS�͵��\�%gP[�`ѕ-����9R���
�ݐ/=l��a^�se-ֈ�W!�Y�#�c��q��%�ʑk�J�MJ�ݙi���R�u��5J���@�.��n�h6ֽW�����sJ��MM�h��n[3�ax����g�<�����5￡m1f��7_z�;���~k��ɼ����+�{���핦�3zJ�Ls�輩չ�/��!�*`ɖ���JJ��J�Hc���@q
W4������z�u��R>����>.���eK݉�ߦ��z-�r'#L��y�����M�'�+n���S�`��}���3�]^3̑\����w8C�n9C�w���M���;)-Ιrߗ6����nM����;HL�d��Y#F��S,[zּ�M�o���;�@zz��V�4�I��u{1���O��(���B3^	m���鞭���}f7�:��DQCRn�h��LZ���g�3��)ۖ����׹�a�J�\�o��H�(�KRq'���L2�d�|&�6ǉx.O��N|B��K�|"����8m�Q|�F����_;'qOD�����n4Ƨ���(�2G��!��/�pʯ�H�^H�k1f��R�q��DD��z���)���'h1(�D�ͩJ�+�)��t�i>��_F�"qM��'�vj�I&�qRF��9��;�;�4�ː�<ԦJ����%QR`h h�����r��
�LI�X)�!9�$��b�Ѳנl��e�n�i�ҠC�|�����S򟉞L��8�w�u���aL�����I9��+��gB�B�)#ӛhe���Л�<A�'%�qGN�ؚk�N��^a��/QJ*E�΀1>��ǰ�d��pS�N���Hi"��G��{�j�iSqRv͹0v����Cqf=�����jjwx���J+��T&Ƚ�(G�I]g4H!I��1&��X�[��L��@Ys����{ܿ�;\k0A�S�IaF�4�5^�w%�\ˑ��q�	����n=6F�M����k�F�!����k�g��j�y��pw:��Y��7F������Fn�4�͕q�V4D%��Q��̑O�t#,�#��{r]��*sFK\F|�-��Z���['T��L���*sd�ҌLU�X�?�EV\�"��W:p���_.�]F���PJXē�&�r���e"$`�+n��F����q����&��7ޫ�5m����C������R�X��+�[��Q���A��儲lZ[�V��bϠ����]l�ϱ�h��=��v �?���>�N��
{���kh�eg�>�, TyPYN��By���/*����ڟ{~N��� �y��<���	��xE�J���$赑�'�%$�d�����3Htμ�"r����IZQv��L)ʮ,A��HI��oF-&%d#4#=^
}�\�e��߳�C��c���hY��z��ԩ�-��>�3D-{0��P�u����_|?T^9#W~;��58jUr����ڄ_J<@gkL:�oB��%��U�}�F�y��z�p�[�{��{�ӆ�iw���������t�����J�]ʁ����b�򨬗șX�H�:17���r,���>�ԥ<�,Õ+����Ri���ğ�o�Q�)���&5d?��d%~��	+.��i��?��?�'�hVc�\�Ƙ!���z��g6����Y������fw�B����6J$�)K ��J)5�-',%�_�Zz�~F����{�ՙ�l��Z��,�ue���bYKa�,�Me�l+c�ك�a����F��l7���v��f���=���}ͮ���6'\�v��y0�Ļ�hޏ��|$O�|���y/�s�C������6�������0?�_���;��	�ʿ�7�-^�0Ūx+�J[ũtV"�e�r����RҔ��e�R��(��|h�Qe��YyZ٥�U(����I��rI��|�|��*�+?)���6ա�V۫�jW5R�Rc�$5EMW�ԩj�:K-Sg���+��ԍ�Vu��[ݧTk�c�i�u����������z]���ֈ�iv�OԂ�NZw-Z��ⵑZ���MҦk�Z�V�����Vi�M�6m��Gۯ���Nh�j�w��O���7��Vga����oikqZ:[",1��{,	�Q�4�x��:Kj<��S��%��h�
ЅF;c��,wM���۪��zH�����e�F���LֵC
��#�®�G��:�.�t��.r�����
�m���J@�UOk�r���l�!E4pu;�OY�����M�d}�8���J����O��,Y��c"��`��_
9H���nϔ�t�4�^:(g��{P'�zB���z�쉕u��W�Y�g���e�tY?,1��z��)ԓ\�d[�$�z��ɔ�1���G˞�Dj!g�����|:^��3� �+dm�ϐu��d���>]x�,Yg�������Y�6��?��)%c|��ϕ�O7�ӛw��0Iի��h��dK�ߡ?�]��v�:Eh�n������	���P��u�k��g�}i]��^�����5�rQGI�"x^w-m6���ƃ�#%摲'�U��ԯo��r������T�1�Y��Mp�}ǚ�{gM���m�G����t��V�RJt�iP=��ߨ���b-ݷE���l2^5�!���/�������7ԟ�6�����-��pm��F�Sj��O��О�Z"��A��	� ���g�\��s�u��J��;]�I�_׳%��r<�q?�s�.b�$W��c9r��gĞ��S\��X����O���Q��xZ�Ru��������-�A�j1KG��Jof��a�����#�L�����^�/e�2A�d�V+ϒPD�Io{�=��ڻ�{�
�`�`2�oN�ړ�{�|�>D��z�zu!_zu��F�y��� ��wNz3�y�7c�m���K�=�-A-z���j�S4a=,�[��T����3E�l�=���"��2b{XY�<�,C�.~�31��T|����{��-��P�cO�Gt��g���@A�`yЂ(��h���J��w��z�~Co�[��1fe�̟�eN֙E�6����(��Ƴ)l+`%���g�٣l{�mfO#Wً��;�N"y�]bW�g�+V˾g?1�+���5o�CyW���A<�'��γ�T��g�2>�?��+�c|#��w��|?�k�1~���/���G��5��o��
Q4Ů�)�J��I�D+��!J�2RIU2�I�t%_)Rʕ���G�U�ze��M٩�Q�+/(��ʫ�y�����rC��ԩL��ު��Vu���5F�ޣ&���4u�:E���%j�:_]�>��Q�P7�O��Խ���zT=��U�R/�W��ԯ�Z�{�'U�ͦ9��Z{-T�Ej}�AZ����h�Z�6U��fie�l�A�am����Q۪��vk���Z�vL;���]���>Ҿо֮k7��b�,�Tڬ�k>����n=��}k�tcu�+;P?�/��$���"<����HQG��"N���1�nV��M�7��H~ˁ��Q0�|��Mj�K�]�)���I�D]�
���?�������NKj�ȟ�io̬���O"�"eGD4P�yG���Mt��\�[�E\�$�	M�e���uf�z���:^��e������z��
�$�_��ߡNV��eO��S�/���hUd�����W/��B�Z�8d�S�ª\m�!����ò�')ɒ탲�-�G~ѿ��MDM�_��IY�n�g��)CA�^帔��Q��GU�J.���z��0���ok��5�T�kZ#��>�;���B��&> ��nqK�U�k�4�E+�iυ�D��KP�uib|�&0pa&�v~V��6i��-0�G`�V�F"�Ӳ-֊UnH��Lp����.-M�|IX;��>]��HߘvV�D���>"�\D��"bq
�4Pg�]�')<Z�$���{��\�%��
i'"x����/���3Ҫ!�*b�h������5"�g�f�p�]NrA�K'���%�RD,Bn���܉��U�o��}CH����#��z��@O�)�<�>�EK~ED�X������a?)b��S�Ej'�OT!���%I�69��!�UD;����?�ߡǦ�K�
���bi��/����m���K�u&GD�
���<]hPAD5=�i�>��7��E���k̻��N̢���`*�yK˘�z��d�M�4|`����X��}IX]��H�ǌa&*��LA$Õg�gH2�gI'�t��L��g
d<Sd��G��	�d@$J>��x��|*���O�����c݉�z�@�:��,��cCX<�RY&�Ħ�|V���\�{��b��&���d{�~��x��^e��;��	�ʾa7�-V��ro���r'��#x���	|O���>��^�����Q��?�7��.�����Q~���o�K�
���k���'�+�bSJk���tU"�>� %VIRR�t%K���*��2e6����ByL٨lUv(��}�A�F9��V^W.(�))_(_+ו��m���jW��@5X�vW��~�5^�����$u������\�!�u��^ݤnSw�{����a����z^}G�@�D��~��Po�uӬ��毵՜Zg-B��h�h	�(-M�M�fhZ�V���k�jk�'�����.m�v@;��Njg���K��3�+�V�^�I�-��fqXZ[�[B-]-��>�A�XK�%ŒnɲL��ZfY�,��=lYay̲Ѳղò۲�r�Rc9f9my�r���#���-�-7-��ĪY�V?k�5�����m�gb�����Z���&���DM���|�+�[EͿh2R��s�v{9�j�ڽ��l�_�|�/�+�ڤ�B���t�~�ɺ/��ظ�Ei'�MǴ��N�����>�����{b�����!!� 2ŀ]�	�P�1�|�U���*� ��+*��PB�����+
2�2�PՇr�Jm�9�r(��R�L0&D���,<�"��ѣ��ivv���{gfw�J�V���ɶ��l�U�;�>��!i�~�r��GI��P��~�����V½�)�^��>Lȶ;���-�y�?�&tG=���+%l���~�^���ބT�����$ģ���=�'a��=���7%{Vo�`��1l9���=��i<�]�$�'
B9�(�M��d3��|�x�P�?��{w�?��v��Bj���>�.����7�7�-$�?l9T�T��@�'|��?�L�Y��2�J�u6��eY.k`[�T����/�}� �������0���gU��^�K�+��*���ɮ��ٷ�Mv�}���}�&�k�>Og��L>��˳�c�'|0��)��/���W���5�v[:!��\ݪn咺]��#j��ʣ�nuOSO�rY=��'Q�\z�e�2��s��������7y�<_����5�
y�\+���F�Yn�[�6�]> ���'���9�C�7�.%��S��J�2D��Rr���$e���*%J��@Y�,U�)+�5�)��e��E١�R�*�)�#���I�r^��\V�)7c,�'1;�ˊ��������&Ħ�f�f2+B�"�!*U����ت�Z�{[��GlB4!�!v"� �����^bGhm�S����إؕ�u<�b,.!І�:g���q��nW�q\����������٢�8�\���cq|b5�Q�؈hD4#Z��6D{�@�0�!N N#�!:��x���bL�"⪉�/�S���l��pΘj.b<bb����%j��E�T�u%b��ZQ7P]�A�f���.�^���A����D=�8��W/���k�o2x��	���Ȁ,Q�0�Gu`,L�t
b����Z�3�z�jX�`-��z�M����}��r�?@��q8g�\B~��ԝ���Pw���Z�6Pç|~a�H5��g�MԦi�d�ᨧ#P{�|5�-��;m����j�wԝ�QkԚ�u��δv��MC�i�7���޴D����n���;u�㨬��tԞ���Qw:�NG��;=W�Oҧ��z�^����E�R}��R_���7��f}��Cߥ�����G�������~Q��_�o��c�aF�1�f�0r���c�1Øi��<�¨2����*c��ި76M�6c����g�7G���)�q��d\1��L�TL�t�Ls�9�|�i�1Ǚ�if�Y`����f��Ĭ1W���Z���h6��f��j�����y�<a�6ϙf�yռavYQ+n��o����!�pk��k��&Yӭ|��*�ʬ�"k���Zi���Y�k����a��Z�Y�#���I�u޺h]��Y7mf�����;�d�G�9�X{�=Şaϴ��R{�]aW���r{���^o�ۛ�&{����c��ۇ��q��}־`_�����[��(��N�3��<�t�8㜉�4'�)p����|��Y��8+��N�S�lt�f��iuڜv�s�9�pN;��ӹ��p�ܨwM�w����w�;��uǻ��錹��BD	��E�u�{]�^��E�uqTu�]�_��E�u�{]�^��E�u�{݃�_��E�u� p��^D\F����Z��^�{���ey��a�/��M�x3��^�W���*�*��[���z�zo���m�vz{�}�~�w�;���z�K��w˗|��}����D���G�c�q�D������l�_�/�k��j�֯�7��~����m~��?��O���s~���_�o�]���x����O�N��i�[��n���(�x��!���7�
��֙�LO��	��(��H~z��(C��F����R�Ҥ�D=�z+�^�Q~��H�#�e��'�n���j��t���!ދ'��{�����{�J�v�l���޽n+e�����	�sOҜT	�U������kz����C�+��d_빵����w��x+�i�	|6�mdأC��>�*?������Mᮓ������9����G�]oe�4��n�}R�y��%U�P~��o(B3rx�I9:�j+dT� �|���$xDJ72k'�b=�US�n�דl����O�����!�Ne�tm'�w&�'����﷙T��p�R�Xz9��R��J�C�l�*�BR�W#!�i��Ie����w^Ee��ʼK�]��q�ָ$�I�M*_I�2�j��R=)?�)"����'c���y�WI��'YG!�F��޵݊��׃�_5u��J�6���`�L�B#>�����q����.��'�j*S���L����O�L5��O������AT� ���x�p~����6@|�L*��J�T��V��<W<�.M��m�;9?E[ݧ���9�x����&��I�%F0�c�$���'�<�牗/!^E���z��M����ۉ?C�Ⳉ�"^N���z�|2�������ksB#vqB�e唥��7e�GS�h�/�zo.��K��xix��
vc�]9��n}'<&l/<�$�o9�r�OQ����T� ����,I�/�"M�̇Lb�����bl/�<��_���l1;®�jz��}v������O:��������$�����%O�s�q�>[�(M�/������ȫ���W#���ȷ"xm�H_�����ק�M{�3����ys�޴����dy2�"�ʵ|�����&���v�^��;�k����jߩ����V�Z����Q�C=�۴� ގ�)S��x-�"��JoK;YEgeS\�����o�W���3��"�2��&��@؈D��%��@����EL�H���;z�ľ&�I���a����b�b-B�q�G��Mb/b�ػ�؇�O߂8?J_�8���b[�Wأ�N�4������2�E�Y������S�a%BV�9�G���$�u`�(���`�Y-�C/jdͬ���6֎~t�c'�iv�u�N����Gy�����y6�Q<����t��y	/��"��/�+���o�|3��w0�@�A��/45��{���z������?@����Kx��&"	%��dk���L�_d��o"!������ģ��W�X��b7`�?����W�$�X⥔.�����y��,�yǑp��H���Dq��)�>�Cќ�"?�q�
�S���H� ޓ�>�elS�{v�@�����0���tL).���B�(.���B�Q\hŅΣ��"�-��"t?�]�X"W��	)$�3k�\6nΜ���e�/�i��+g�����%� 3f�⊅s*��E:��e嬲J�\B-гx����}��4J�;R�;]�bA��U��ğ�ư�lJ"�t~��B,!�ŉ�ŞN���bp#=;�><J��ڠ~W�:)�WI�T�GH�E����|=�J&$��t���v ���wþ�$��Ⓝ�䷥�������ے��K?�[�����S}��X���}�G��Nʦ�"���h�El4<����<S���E�3�sx��`.������_�W�5x���߄7�;�=x~��m�����k�����Q�b�X���;���P���=�F�W኶/E�<�ӆ��Eb3��0� _�/�_�_�X��U�k��|�ހo����}�l������G����~��
T�� G��` �1<!�5Z�1 Z-A�,�������X`F���Q��,#�K��cL�|(�"(��P	U�j`9��հ�A�C4Bl���S��^U;�K�u�2ġ�`�]�	Y��򧒃�,�3h=h���$�J�'	&a�ߥQO�D��3����`��@+�O�=�c:��μKg�ՒIEQ4"^�}Q=O6*lk*� ��x�]˕p��hõ�R,{��a��?��yG�n�Wq��C��8��?�?
endstream
endobj
20 0 obj
<<
/Filter /FlateDecode
/Length 467
>>
stream
H�\�݊�@�_�\�^��	!kF�����} ���0Q阋���]��a�D��ҪN��p����a�N~��0��ߧG�<��uIH�n�*�w�v�"�O���o��2�nGů�x_^��t�_��z��J/�Sԧ�<��*�������o����y*������ay�FϿ���'���1�������ve�*�5�ȏ��6�Η�i��֛,ӭ�C9��P�j�@ᡀ]�����A�{
��`
a�`��`��`��`�`�`��`��`��`��j�G� B��sM�Њ�Ԛ�Ԇ��0H�Ўc�[�N��>pX��@��@��@��@��͆�4{^�4�������U��Ͱ�jkx1�a�C6�B���״xh@�済d�8�p��].�[B8́��!\Ɗ�.�D$�Mc��k�������B�t���^gy��y3O��J�� S�t
endstream
endobj
25 0 obj
<<
/Filter /FlateDecode
/Length 14523
/Length1 34888
/Type /Stream
>>
stream
x��}|Tյ��g�s&���+�+�$IHe��< Ɍ3^��O�(-�"���H_�����km�^h����z-�j��49���>g&���m��������^g���^{���^{�9�㌱� *sW�>s�s�6g;`vaQ�wzMc��ͮ(���s�|����^9�ja�g�	3v�P�˫��ޑ��m���h����ퟶ瑧��"�nu��X�ã�mn��7�\5a�J�2Π��9�X�����g>�Lc,�Ř�T���3ٯЗ���D���{p?��%��Ǐ��n������W羶�53��6�?kq��'�j�~3�Z�-ޫ�8~���m���7��1~:��^��gl�^�wF�J�������ʤa��}^{v��ȵ�����o��֪��9Ź��J{�yF����Q	c�f#$�$@2�#
�!��EC}Ey�A�x���Ͱ��7�^�NG��UEQ?aY�W���B#�cE}����+�S�T����?\����w����F�*3��}�����l��_�'�u����c�3�*v5{��V϶��-l��gx�����LG�l���gGX�Y��El[�� ߄^K�J6����A�T���_�+�v�]�v�X-zoE:��J�kQ��A���eh?�M���+��'���8O�8`�1R�kX�,���Q����A�|��Tޓ=���t�w&)��頝��!�ք�B
+Ł���{gJD�H˭v��2DR�)�4�MǨWD3��o�2Q��@-6�~�	fH�u��3,3��!��19�[62���6�v#�Fs!$�	spk��M���K17����/�'�bH>����h62��,��i;sK97�f��,X�!磗��
�F��R�lYO��7Inj1�����h�,K!�@� �K@j��u[ �1Y	 ��E��e�YbІ��CQ���W�m`)}�}|�����Q(_ʾ�]	<���$Уu���Ѱl��K&�^���f�'|V�:@�jdf��T�Ao-�v��ϊ�r�A7�êoe)��S��2�dw"נ.��Aߔ�`	k�b����(܌���ٿb�(M����U�;�r�j��e��4zj��k!Y#�8چ4R�*��-`s����3��S	��|!R�c�p�O��H����9�s����P�#y�߃Du9|3�v��7�H�y>��s9G���Ķ���/�%>G��cF,�#A7����\_�3����2$�W�{���">���U�X���w;�v�� Z/g����O��S�,z��s������� �Ϡ�������m�xc��g���u���fr�z�(������[1�a���ץ�[1ӵ��8��c��>��=�Ld�(� ��➼��Chu^��V��ɵ��R��V��d�Z�<�gM,��21��'���,�ð�'H
d���Jk|x[�9�a����w�c��z��/Y*0m� ��>$�����6�6�������)���!���5�3V��G�w�eh�Ⱦ/�<9IqPr��Z[t���{z���HC�-���;�Vx�!����A9�}mƢD�i�"�0�O;�޶��*s������\�^v�������D蒟�m��h��*�AM�C�l�/�;	c�іv�Z�\?�h�W�n#����2�"�f>fq�l33�x?(��AXY;y
ی<BF�g�R>�������@��X��1Fx�������q���/��i��S�F��,V�t$
���%�N�������Rd�߀#����O٧��f�g��J??��	��.��f`�8�%���G|�(�L>��"M��y3�5�Q�i=�K�G�6��?&Y���1��h��@7�&�y��'�Om�>g���l"�i�6 U#�OD~�̃��ȃ@y"جDZվ��c���M<>|2�W�e����)(5B[�?tH���ex�[��O�/1샵��ZX�R�:�Ԃ����`���^�1㉲v$�h4;�N�L���F�i��@���eυ����H�q�? i(R|n���F9r&���,\�,DMV˧�ʖ��z�ͅ'�E�p~�pDr�Hke/�����j�K_�g÷瀇L��(���HT�=�FVG�"eD;�dl�V�f�(*���R�-��S�L딼 eM�䯋��QM�M����-�).���(zf�����.9V��؄"��LcS<����ʓ����;;;�4�2'��Ù�	�c����pJ8�����:;&I�ގ��w�w۷�o���P��XU���{3nȾ�?���3�c����2Խ��3��4�`�d^���~O���r]R�%�\f�1�77HމW��<QR.��^�7���|��;<��E�!6��B��/H����4�����v�]�ԑ��o��9�|�@gQlG�k�����lv�������S[���
|���Fg�1�2�Z2
[�cmm�i���6�ns�5K�%�R��=�3#�߇�_����,�V� ���$JǐJP7��p_S?�L��h���q�4���{�pyގ�pb�\i�}Q�ft���Jk��g[P�&��\��\{��!�8#��h��e>��䁀�pM��aF�N��� Mg%1u�r��JS�O�[R~�K�LXӓ����Z�WC�0���.t)o`� m��1���,���
��ly�J�ZS�e���]&O�:��q�uhWîb�xX�%2=j�3qJ?b�m��8��͟,���Fv֯I���-@�ނ"̲o�ٽ��ʱ���H���~���LY)�z���g�?ԄͰم�ץ����<��Dk����zPF�ٰS��j����S�=��<�':b�h_�s���NL׻Od����OJ<c���8�Z�R�Zmi���@�� q��R&�c��Y��NQ�*?�G�ʟ*��}��f)�m�d�;����t֊�礒Οǚ�{U�	���js��H����R���I�׵|md���MJ���8n$dk�t�|�4Y�6|R-���ɧ~��;$\)�뎋^�G��Tu>�O��NeJ]�[��5��26}I�Ys"���iH�Û�fI�n'�{��G��}n�.C��)������nA�-�>�h�������x�`P���G�܅��߰�~���:;�5U�~�}b"�L`���B��)�]��i|�g�;�o%��g���md���:q��� "����B�6&��P���@!
�2g�1X�9�+�݌��c':lGD7��M81��^5R�~d���N��4�9g�K�e��1�Y�Ӂف��6o�9.�O���aׂ�q�v���}4Z��l#�_F��М
��+y�A�Cqw	�� �'i蓋Xyv�\�h��DM�Ov�ҟ�������������]"�%��|�}�E��%R_�7��B2��Z8	�
�	�/�"Mļҩ�F�.��jÌ���ɒV�/R�2���-�d�û(��0������*�d�j~	��}����yl�&p�R��g�|�ߵ�fmaE5/��l��"��d�|6�)��g�f�!�R6�+7����Z-�ڀ]����m����r�:�+���┻�2΢�?�^{�߇t2�����ӕ�C�#�'t��(c�:'y���o�y�P�~o(����.��Ogn���W{����a��|�W�C�ǐ�����~;z�ê%���=y��e��,����Y�[~�W���/���^n�)|3f��O�J��!������;�wa/>��c�>������$g�w	Ǜ������>��/'�����J�@�gh�>J>����/l�*��a����'������JDx�p����/�*�xn:�W�cH�yb�}�6O�v&^g!���,F�YYyr��I�p>�X�r;S�^�\�<	�J;S��3�
�y!�����/�����X��u�Ξ�g?Y�bI�-K��1�4BRM>o��hi��/d�~��5U(�e��+�J<��Ը�_2xLv�[W��u�U��u4��Q�kKk�aq��aC������dϫ�q~��ЦZ�����h��
ezX�%+��]�%�6d�m��ic�Qec^�)�|R<���Y���㳵#O��g��rţ��#��a�8�]<t����*q��8�K<h���C;pV�k���-�~S�Z}`��-⁍�ei���}yꏲ�^Sܟ+����;[�����V��a�v�l��|�����U��b�)�9+v��7Ŏ��_�����.Sl3�wMq�)�z������jw��۷$k���-��;��wr�m��u�ڭ��|�rm�b�F����i�,��77ݘ���Wܘ$n�.�7�&�۔+6^�K�����n<�*q5(^�+֣��\�.]�b�G�1�jS��=�`�*G���G���֖'�VS�4/�Z�-��aZ�rќ��Z%V�f哢)/<L4�O�G4�����>Cx���u��5�{�Xa�+<b���2S\�*��%czjK�DM�X�zj�M�(W,4Eu�S�NUNQ� M��.T$k�DE�(7E�|�V�]���RS�3�ܒ^�����sV�>+�7���^Z�Q�K�J���\13E\:#Q��3�;��b�SL��G��]L��Ԧ�S7�S�bJ�:yR�6y���&���ҵ��Ą�ڄt1>U�^���z�%��$]������+c�EP9bLv�6��sT�ˋW�G'i�)"���p7zT�6:I�>ʟ��(=A�(F���#�Ib�<�54]�*��2l�
�MCRE�T-3WvM��.�]Ġ��ڠ~"�SD���b@��߯��Z�j��)Z�^���S߸$�o��K<-V�SE�y"�Ҷ�ޓE�dыgh�Ί��"%9WK9+�Q��+�k��"w�5�����3I32�3I$ �0��$gI耄C8H�xU��5=A�Gy�c�/�����U��B(=4�(8h��z
~�{n����_�a���>�x>�ⷳ#�u�t���e�j�;�G�ǖ��3�2��2�F�+�B�xD˵�3���6BI5�ITC���Ml�xQ� k>W�*/*[���D^����I�)�O��0`�����F?�����<�Oe��E�����^�8�{�΂*�^gϱ��k������|]��]�UlD��z�c$�l�	��O�D��s�1�^٩<����j�8�,S�Vv���� {WO�x7��8�*jO������3�����D�v+��8����r)�J�\l�8�1�T�ݱGO�c�i��;�p�ƩBa��v�Qۋ�����1��qZ�����O���%�8y��^)�S�Nܨ������{s�#�̗}$h|"�O���S��8��j\�N� �g��;��%�I��^�\���hʈ�v�?T���,'�_�M̗�=6�d|���5�`�����O�S�>y�d�N��ȇ�XJ2���'%��Tz���;i�:�x�B�U�Y>��,�UX��tϏ~���C��;�Z���1t�y�8�w����bҪ�bj�c)lD^o��pr������=2XR|fO0�~2e*>�����a̔�!|�dg$�+�}�!�V>����<������q���	��f���@��A��� ��̸�?��E\�M)����ָ@���郝3h���ǣ�0O�J�95e긼���Ab��U�I<III���/�)C&N9GSz�Ԕh�a�m�;�q~��P���V��w��s
y"x���d��Ia�Ǚ?�X�a��f����8��:�r�!y)���'^�;tEM�c	F����sIM��O�JS���b��>��>R}��f{�x���XiD�}нt5��g�eJ�ڟ�!>�`�G'Ǎ�d��Õ5��k�S�E�w5������8�Z�>L�H���&��-ϙ�P�������(�8���R��8������CT�H�~�HV��rI�#[�9_�W���_��T.U.��,�e��㡄�9~����]|�+&�|<E\&n��mb��%~c������{���Ş����#qO��[Ζ�;�P]�$K��6N������|pʐ1D�Y�W<�0�5w��^��*e�������r�߫�~����`KN�3�K�Ä�Z{��������R	��$��a�i��r��e$.�4^��xU����z�Wy��W���0��~��g��_�P��S�����Zs�y���o�l���p�ϛ��[�:�OLJN����5�jBƦ����~	��}=�zk����R����C��JN(2G$�����j�\�4]rn��}Y��s��	C�G��wj� ��{���3���dpH:qB�pn����6�����U���{���K߻�����emE��uᓻ����Yŋ*f.�d\�[�>xw�~IueݒYށdoKao0?˃�_��d�����t,��H��)��o͛ԁȯq�4�LiT_1���8��S��t��x���W`׿;v��MK������ 6)o 뗨��~����q��[yH�QY�����9P�r�\yr��E��j�቉�)S����xj��(K��Cͷ�~�����b�Vsw�W��^ye�xF����}�Z>���|�r3i�ѣ{����Z���R�ȼ��T��REcʭƝ	=�Ә�7tq�X''��X���q$���Q�L�nܦ�˿�����6��53�������Yͭ��C+���_f4���6v���{�2�V���gJ���(Ϟ7�Ib����t1]L��t1]L��t1]L��t1]L��t1]L��t1]LSg��z�xb��/�d����,wVYa*��e�zG�jLYc�e��b�2=��.;�@��.�����i��F'��x�KXe�9s9G�e��9��e�FE�jLYc��*���,g�N�t~�.;�4�v�G�,��]Nd��Gg���M�!׈����q�ƻj׹
�B�P��n�v�����]��*�����^ONB�w�{Q��������������o�mn�sy|-��H�*wk�5���s��=���`��Օ�3~�Հ�zU�}�}�.&C!���c=��n�	��u�z_������]Ӵ�ilS�ǻ6���[�T�mz�eo�����z]��fߚ�9�o!ANBBgg0�vY��zKs�OB�?�aW�����+p{�-��*���;���
o��)(��֍ހc5ܭ!�'�U������lW��r��s�1��A���R��e��kO������Gsjj�fKӮ�R%�#A��r���&7ƃ��Z��!w���oj��GE��U����3GJN^��i��J2�&�T��J�t��,�5�y��5M�F_[̴4�Q���J�m�=���j�J����c�Ȧ1������M`�������I�![ur�5���s;�4ԷZ1�Wv��\A_�+�V��["���f�$	T�k�4��i		ըr��V{��I�F��a��f��iV�+��P�^[k`F��"��vp�����
��{��(�b�km�{�o�y������!�
 ��x���h}�૭��y����V�FC�:c�:����@$H="���dY��R��9�@7"v�/��bk�:WSS�H/��K��B��IsY"^؝�`�/�	�2�k1�ƎT�2i�fJ�avl�^���j恄X�k�2�]ªq��~,1wm��*,�A���4�C�Fw��]���:-��j�������W2-	/4�A�e�l9u4QnW3y��HC��n���a-��G�Ƿ7�.C�i�Eos=15��U\^V�*/�^�_Y�*�rUT�/*),*te�W�>3۵��zN��jZT�U/q���˖�敔f��j**���\啮���%E����*]XXR6�U�~e�ծҒ�%� Z].�ڤJ�������Ysp�_PRZR�$�U\R]F4�A4�U�_Y]2kai~��baeEyUh�lYIYq%F)�_!@hVyŒʒ�s��ѩ�lWue~a����y��a9D�t�&9�4\E��s՜��RWAIuUueQ�|jKڙ]V>�t���0�����UPQ�J�,� ʬ����ٮ�������:�f�8����ʊ*�K�]UE�J� =�Tͪ�-�{h�T�;����h�B �.2&dN����,ə�������(+�K���]��%U�Bqe9إ�D�q!�I�Wf�KsD�s����-`aQ~)V紅u����Cd���ܣt���̖Vk9���V,\'��g�,��X�sqі�m�_r�n�F������ɕ`}�ș�i
ʕ�m��g�{Aw3C�h+�Kw3��lv]P��hB�5������l�i��쭪�4Jw�ޠ;U�jo���~&9ijE�b�.�W��!W�$����r\	l�!�^���5�F�.6�ձ���qH�Q�E+@�"�W�h&�֊�9(����b�QZAy��Ջ>�=h��
QZ	
�XZԡ�TdK�D�*��~�
�f����~[Ђ�ө�T��|�jE&�}��A� �~>I5|�g��P�����u�zYoI�5A҆��4�_�=v��h��v>\��+���9�%j!�^�V!��RQߵ�����R)�Wr�e�1cG���s������7�a��r��{� G���|#[w����� ���?�h��	v}��M�]��-g�Ejup>��7�B�UHz-�Z��Z�e�ז�A��*��#���Zot4k�-�˖|�$�����^�>P�3�$����t�fHr�uE�ѪNZ�ߦ�@�-ޛ��4�Vf��dʙs˵@נ�}ܶ|���*[$�����^w�l��(��#�� �CX��ӈ�:!�ЇQ�$���x�!ik��Ȑ�����#d�k���I*�N�Hh�"dk�E�b%��t�J��6���١r����\w�� zg��Q9�J/咔��`�n���u�/,uDs���E��Y]�Dk�>Z����P/=l�-�7fD��4F����ׂz!Q(�&֎�m/��:9�Gr�ds:M��j��|�'=C����N��	h�	٫!إmd����b����n{�j�~;bk�6,O��|����E^���٦6�$����.��P_�ɺ(�-r�5ɵ�h�{��z���-_X�9�VٿhK_m���"y$�4_�1�h�/��]8)�C��z,ۍ��]?�o�)��y�X�[���8�0']�뮗��m�{���t��=�W��҅n�Zfd�t�E����v��5R*��y�}13*w��>��f�X��vJ��3�r��bxm��Cd&V���<��,d�5�ڏd�bn�Y����o�|��(=�K^�6�^iQ_o/�t���T�fG���ʼ`���e��5��e�-Id�EVE��$`��J�/-z`�=c־hE�����륪��H��룚����8�w4N9��bē���^v�/�.��K}!Ӽ���ϔ�q1�D�\�t�eӨ$�K�!�.yOw�о��o��cɗ�P�JI{>������
i!�<�Q4j�W&_���K^,N����+W%r�g�qW	�s��|�.���l�)*�E�,�9͗:"�Ds8*�w�]�k�|II��G��m�����,E�k&,�f�Z����lz5��F��[fK	I�BٟF�'�g��,S��J��K��|%qQ�H~zI�K�_L���|ЏЍ��lIa~ԎJ�������H�,������YR_4o�y�)_j�꼒D�u���YGd��R�"��Rٺ
z,B��(Ʋ�)�,[�M��-�(���,)#���Zd�T��]W)�B�wJa�@�g��s���ٝ��rie�je�\�E�U��모����os�0��"�ж��(g]�YG�v��wX�"cw��BiO�6�UQm|3]�wa_���k_#��u玍;����3�u���H��³eۖn�:������3Olw��+rJ�b���7}X��:�F��[�`0�X��/�����{�ul�-b�{A9�%Y�ݣ;-+�t�h�F�G�ڡ���r��FY#�!;2!��춄_��T�v���9���M����3�L�$5L�d�M7�"�N�����Z��z���i�{J:h���cϸ����`�!���m��{s����o�Jd�~���Pna\٬|���N��Q~��n�j��k�[�P7�������(�����k�{(����q�Ώ����q�q�a�(S���H*��AEc&�C�3��V�,w�]��խ4���*V����زfw�JS�4a��VI���xUe�8n�pnYaX\I�|�0O�R	痗��2}?�&Tͫ"(1�t�&�'a��9-�ZVQ���U�/Ka:�����9���,�`C1����R� ]R�c_[ї�G���p~�u�ѺO�#��,����}�S��� 3�!����zWo�p��>|�,�8��S���i�7HG���M�
�:u�z��!��T�~�J] �\])ˍhy3�ٳ��zB�I�i)���h� ����Ō��(fm�1Px>|�6T�ʮ��(��{�M^��(&5��	5���(\y!L�,KdR�k�M��9�s[W(���%��o�����)?�O�
St�Pz*�J�2T��S&)3�e�R�T+K�J�Ҭ��ʵʍ�mʝ�ve��GٯRS�P�V~���������|�|�|�|��EĉD�*�	���"WL3E��+*�"�LԊF�*Bb��(n[�6�C�{�qXO�g���%qB�%����KqF���&��j�:@�TG�9�u�����j�Z�^�zԕ�_]�U}=�����N�^u�zP}D=�S����*C}[�@�T=��V�jL�5C멥k�Pm�6N����
�9Z�V�-�Vh�Z���j�j7j�iwj۵]�m�vH{L{B{Z������������������֮+z������t���g��}�^���+�E�2�Vo�[���^ߨ߬oѷ�;���^��~X?�?�?�?���������?�O�_�gtӡ:Ɏ4� G�c�#�1�1͑�(v�:*5�+�J�߱�q����i�fZCJ�Y
�(mu�	kWf�k k�k�pF,P�t<&{�V���6`v���f*`��N�� Ie�1�#W�O��&O�τ�\h&�ˀy�\�6�A�U0��|8¼P���[���X����Ą�P����u��+�E1[h\ebx.�	��w���L?`K�5I��ZC�uLl�`�a���xe~Ga���֑,Gɐ���$�R	/��4�K�	S"�b����j9A�y�� ?Ƭ��y��e�"������Z�Z	C4�|w�_�������_���4W�Y;@�Ǵ?ޑ-g�I��93��2��Ae���p`��PB�{�\���솯{"��,î0�19���+%<ɜ�M� |��9���t�\n���;�������*@��@s-a�9���	�?�Z�G�kp�J�&�[�B�ic*=� S�nc�|I�;������� ��w�/?/|��O��u ���$��~_b���k�/e�K�x�m�:j�
��A`n��%�V���%1�a���(t� Mw����ӌ���2Γ���%r]���͑l�������c�҂ްpɢ,0grs,�_z��T�tȱ�5\.�Icr�{M��o;~��f����RW?
��< 4�rW��6�f5Y��$=C�(K�r�<�B�4I�0)��y�:�E�y�]�kΔ��mI��<A]�.F�u��C�E}�e"�t���#����F63�l�1��Z���I��q��;�_�����F6�t��np,���(ꆩs�톙7��]�?�aLgd�}|��߮WoPoToB�N�Ko��w�һW��)g2뭴����+�Hr�E~K�Y�Xo�#>��J�v�F;����K O��g�s�oW%NITR�~�K�R��\e�2S)T�*�"e�R�4*�JHY�lTnV�(۔�ne�r@9�Q�R�U�W^RN(o)�)+'�/�3�)T� �E� 2��#&�i"O�RQ)j��#V
�X-�׋��q��)���A�8*����W�e�x[| >��iqVe��jO5]�P����q�$u�Z��Q��ju��B�W�Հ��s�z�z��]ݥ�Q������'ԧ՟�/���o�������_�횢�i�Z��OsiYZ���M�fj��\�B[�-�j�F�Ui뵍���m��Cۭ��h��#�Sڳ���K�	�-�=�c���vF3uUOГ�4}�����s�	�4=O/�K�J�F�B��+u��Z�F�^߬ߡ߭�������G���1���+�e��m��S��~Z?�`�a8z:����Q�q�I���G��ڱԱ�Q�hvk�:nt��ӱ�A�#����8��kߡ���s�+#ee���%�v�~*�>_j� �����U�k��~v+�� ���
���
��1�x��X|�J�-G���)�#Z/��N��
�$�a�Pt��S_e�N�(�寒��o��V%K��g�!��I����#�1K�$����*�u�?*���3�����k��!�J�J�s�F����X��1�&	�$����K8M�	WHx�J�T�J�2��4��;IZyc���5:IUk�2][M�VÙF����V��������� ��AQM��Z��N�i���S�~��=R��y�O`��U��j��]M��o�Z�G��(��ZAx�"����Q�qu��S�\��'�q��L��w��"�/H��C�����j���3�O%�4AGI�n�@��Y�QT6+�4V��w���GVܓ�K�(vZ*u����$j�a�ى2Y�'-i4��:�ܭ?*m�(��v5��Rr��j��A[L�J��(u<QP�$!�z_i�|@��? {槴p�JQ�z�����^�k��6�v�I�u��+�#Y�6���~�QT�.���F�B����ڇ֚�ߪ���H �_����U��8x�Ng�QN�0G��KEk9���V�E|ʙ]�RL��XG<C�����n�{}�tH�5�	Q�o�����G�Ov�V7�P�w�������XI n��l��Hv�#��oj	?J�F��B�R9S<��W��lI�uZ���R�"�!�sW�	�<([��p���d����Ng�[�3RK��� yI�L_�(� ����2O����>��Ho�G���K�tDR8��&�+�Ij��!gJ�/=�C_��i�i�ɳ�gu�Gt:��=��ˉ��pQ>%���/ Rp�Ԓh5TFPeu����d�θ�(`�"�Q��8�3G}�?e�/��Q�C�q-3��x2O���5���	|��ż�W�~����W�k��|3����w�{�>~�?�c�8������_���7�,Ҷ_��G%�$�z	wK�3�M�9�skυ��E���WW���<Sn�)Ƕ�)an,���o�~},Wߦ,)��.�M�f$~������|6|{I�>�O�$��e1\���)�Y���	PQ<�	��@���`51��b���|Y(GN�k�\�%�o�o�\*��<����r�A��i�����L����4�^��&�TޛM���M���<���_a3���cv)���fb������,+PpFf�p�8�
>�H����u�V.�w3��O�a�-�-�ɱձ��tls��V!&��Z������y�� �;��18;fA�c��Y��u�l��?��u��n�t���*=Yo�[�\�L�#ҊB^���f�-����
�y/����G��B~�y��I��!N����v��>Ȋ�=?�����z����ٶA�ݐ� �9Y��/��-������s����?���(�@�����U:.���G˯j��⿮���]9v��Wp}T}Q>�R��?&��q���=�
���9=���in�4g������LO�� o��WHx�������p��`�Y�{��˳�\���X>k���k��昧��O5�)�C>����Q;��IƊ�sV~��UUU ��/�O k����F>���O k��Z��F>���>��Q�,gz��d|�;�eS<�Mlf}S��6�6��\ ܬ��W��I����ib�j��"�)����G>[$�v��Cj�}�i��c_K�SO�}���u�K�/��o_�Xc)��~J��|C>�'�	Lq~@O�Q�+��??�ԙF�Q`��\�Ԩ0*�E�R�
�֨7��F��j���z�Z�z�f�6�c����i�6����A���K���Ϝ_9O	�n$=�t#�i��c�1�Ȥ�o�� Zgj {`_-1�h��+�z�1�(3��c����~#d�5�167��-Ɲ���c�q����o�0;۝���:O:�8?7#�H6Rf0\F�n�ũ�3�
�
X�
���	8�(���i��^���O�~�|�6�U�b�r�J���Ac�q�q�q�q��c�q��/�=�������Cο;������_�2���H2z9�Fc�1����Y���T� �'L1���Q��`�]�CP����8��R��QSh<
�g<83ZsD�<&k�5�T�I˕߄���r燀��bKP2�0�0��q X��<b[1>/\�����ڳ#������<��
endstream
endobj
28 0 obj
<<
/Filter /FlateDecode
/Length 263
>>
stream
H�\��j�0�_E��P�:�F!JF!�}�l��JfXl�8���l+t0�-~��B�Y�=wF`�����(��]�Dp����a���Y8`Q�oK��3�����K���� ��+��Lp�j������h��i@���*f�e�NŸ�1j�2>7��3��6���	�^�	�>��@}��4�_�B�a��§l��$S��'���JDN�]�nD�,89�YQ͂��,)����>R�i��%���8�y<��޿�Y�T��
0 ���q
endstream
endobj
29 0 obj
<<
/Filter /FlateDecode
/Length 759
>>
stream
H��WK��0��W�\X��-A	4f��[��Rzh�-�{���Cg$%�Ҍ�Cp<��o>}��>��v�<$˫�;)��r���ׁ���A��KZ���5�_��^ z�q��8���e l�6r���k���PO ��7���iޏ�(�2�a�(T"����I-%�N��nj/Z���m��\Ao(�$Gb�'Qc�i6����ƿ͟ON�TPp��H&�O�I���_����f.�x�
�9�F���g�Ll����y�b��Lx����C�����&�.0�91�qI^��w�{1ڌ��(aݒ�������*]T��y�圀�B��
�!ɞ8}(!���ݩ��lv_�x�|��H�e:�L�p���a"��[����bo�P[l��n���bJ#�7ru�CF�e��^ ����)�rZ�6�$�I�0�$ L��WIЭZ�U�h���A���q@�~:��6��6.c����+4���/�*���w�_^��C S�f��
��˰
�+��
�k�.zJ��:�������e:����?9��Y�)��@$�	���ψ��7���� Y7�|{6�D����m"�?�M�P��(&�Z��b�w������iA��� 7�Y�����n�ڻ�Gz���Y-�wH��"�(�}�|n���iX�i85��Y��t^Z��9ĥ�K��v��p���9U�5�N�A
�S�f#��=;سI5����=������w���n�[����h�'� �d��
endstream
endobj
30 0 obj
<<
/Filter /FlateDecode
/Length 541
>>
stream
H��KK�@���+�z�W&	H��v�N�Ną�"v���W;5�q�ם��4��39N�F� m�.�~�*�/ĝ����x,¨Ӎs\������w�����=N"�x=�{bk�8�ĕ�jX�ob3NK-�tu3��à����,�ɴ*5�ʩ���Z�-읕��mI	FBϮ BK�� �Dj�AKJ�Z�.!Q�\�=X�/!RK)�2�͘�u.8	�
"����8��͘�u{B�`�o�D-�87�� g��u.�f��X
W��Gs"��䱚T ��G9v�\��4��Uˇ���8�tX�.	̩���2JKf�]�߃��0�Qs�֏���y��7Q�N�q�_��p�j<���8�W�+m����Yc-�`�1I�X�R���v��7������`I�H��xdz��ђ�f��Ǟ�%�e9�?LJ�o�ѓs/c�(C�9���}�Y3��R<c�&�g���59.1[��G���O��YC�V6n�L�C�T�h��@�2g[DD�į4+gJWȅ�����W5���c@�%� j���
endstream
endobj
31 0 obj
<<
/Filter /FlateDecode
/Length 661
>>
stream
H��V=�1��Wl�t��%����C�!
��Kq��flo����I|�V�x'�o���Rx;J���	gFg��0��ე�q3���e���C�<��Ҍ?�����k����������,�<���=<��^��Ŕ �q!��?��r��l�p�������X��n�'��T �ꀥ�X���-�%	��%����sH�U�7(`�����0�x�)c�E�Z4�-���w8����,l&���c��o��_�StRtI��y�/����9![g&)��&Z:�w��"h7�O'��F�j��i/%�b� .|�����]��X�A>2�YE�%�Bd��,�R�%K~8�8~4C �:�A� s��.:n��+o�`aCZ��,<���SZ(�C!���B�F��!�g��s���s.u��Am�JM�ص
/Z4�6�*�s�`˜k��$�Ե�8�+z�i�@��8PעEhV���u��Qz�=Ec ��̆I�y���̒1t���":ɺ�U�LI�Z\(���;*.3yY���V^ˏ���[D�?��ne^��X.�t��D­��e#�(���MA�nmPt�0�,�?�kj����*����	���X�7ˠ�N(����J7�[��}^�U�D˨+�z���L��}����t�
0 ��Y
endstream
endobj
32 0 obj
<<
/Filter /FlateDecode
/Length 579
>>
stream
H���M��0���>v��H���a{��[�Ж�9���P}9xv5��LFʇ_?zg2����0�A��S��v��?N�����ߟT���?e44��>�~�����ӽ!�:�&��ܠ˝��Y=��>�Է�Z<<EH�������z�,4!�27�-`er�˼�j��
c�>�?8j��[�P40��L`F�ջ�	�Ñy�X�����8�VpާˮCj�|X��_�q!�Ʈa�XV&�{�蟗�p�;̯}����h�♇��� �*����B��q�u+D�%N|f!��0TU��h��|�Pew�0���M�8x��.Qew:l�[!�,qb�!&x@4��NReƍ��fS�M��|�.�Ʊ����|�,����Ɓگ)Fްyklقŭi�Ě#k�K�|�.���X�w�$����t-�H��!)e����#�(�<����q��<rdB]=A���6��e�]V�&^
�]d��J	��4�\�v����<�9�I��	�}��ǉ?��)?�Ż�@��w������[{�&K �I��B{s6+�$L{[��H%mL�=3� jm��
endstream
endobj
33 0 obj
<<
/Filter /FlateDecode
/Length 603
>>
stream
H��=��0�{�
ׁ#id�pd�HpR�n���/n�aG�z��+��xW6˫��hF�{ 0�/�<�7���sF
���^K�og�:���C�������5���t���.>���G�����Ngq����(��!��V�8�İj��o�R����/�	�:�Q&<�:}Z�uJ�}ς�%`���ۈ��41����x��a��aV��6Z�Á�%�:�4(i6�G��C����E?>�>_X�z���j#v&�,[i� k��(�&�$H����Xm��<��b�}�=.��|a�#kUV}@��le�z�j#~&$�������<C3벘ቮ�(�l ��N�k���v��U��y��5�m}=xqTrym�ojdߒ*�����=Wտ��B��A��<fki��1~zbo�E3 ���>]�D�:PK�7��:��[$�K�Դ]�}��I��%���B��=A� 4� ���D�A=s�&���i�-�Sܽ҂(x�ս�oqR�	h���,|>:	`���K\ho8z��0�q|��s��_�C��)�H��υ�#��<7����*��4����8��'�Y���+��T,dT�.� *���
endstream
endobj
34 0 obj
<<
/Filter /FlateDecode
/Length 604
>>
stream
H��M��0���>Vh�m(�t��[���S�-�9����3���ģ��P(!�b�W�^�F# _�5��$���R�T�s��&>��$�n����J��%���x��2��O�<���>,��T{����I@'�E��Њ� G�ChCω"���P~�ʚ-���>�CO�Q*� ;?�2}�ƍ��ж[6k^�-�m�7:i+��:�8y��.k����ڥ�H�����d���G�!}�YR�9ޓj������.Ѵʲm�/���"۔��ԭ;D�ms�FY1�o&ʃ��T��,�e٘���K뎬u�W�~Y�m�����3Dj�O�y�r�\(���W�]����Qj���ur��71�!�.�=�m; HFR_f�9 v�x��
�4>��V�|��;U����>�T���=y�k+դZ"�<���ӟ!�6�@������z��;o�(vV�J�\k�"�hM���fH�%�vo]��3$��9�9O{���<W8ū�DU ������qrP-��,|�~
��;϶��MG��T�΍+�t����U�b_�n)o0�����9�1ķV�Y�ѿ��n��̏+��Ž�Kë  ���
endstream
endobj
35 0 obj
<<
/Filter /FlateDecode
/Length 601
>>
stream
H��M�1���>��C�x�����JO���͡���J��oF^'q
�2$�L<�K�,ki�� ���M|���j�R�EQH�'5����Z����Jk#�q�/�G�_�w���A++�	��׽0����uًIE��Sn@��HY����-?��t�C�]CX�BL����)oEn51��r�M*5[�r�~W�,=`�gՠ�7Y�<����������1v38e��\ +sy�&�\�8e������}�f�Qp�Knu�{Rm� ���6$�j�"�iT�@dپ,`�R��(����|��2Q������,e�!ncVVѯL��5�����v�oBu���B�ȭ��a��V>�{��*=��h^)Ӝ���E�M�7�y��9�m; P�@�W���d0��D�[���/���V�hiC�]���y�K+դZ!�<B�6�!��ځ6�0f��8�$�+�q��q�f�b�5��R�d�^Ӕ��`��Z!��ځj8C�� ���4`m1p[�/7Ҍx���K��9���pi�j�S�i���Sm0�6�ח/�ֆ��xĊe}v���t�g���eR�9���#� M�R
endstream
endobj
36 0 obj
<<
/Filter /FlateDecode
/Length 564
>>
stream
H��?O�0�w��H���	u ����1!B� ��W��i}!4ɀ��6�6}����%A����D�ZV5&h��y�
����U�.[a<���&W���&~����˅x�����u���+�2�FeoH�ۊ+Dԫ�]��S���!$�]Q��2$�A���Iv�F�u<D\,�E��cd��c�w�� q��7
WO�}���]r�5Yv�5a��Z"(�#8�Z$˖r�Ax��)�Si}ڎ�C�g7�:E��f�E�I�6[�H���F�d���L�o��=��c(M����!��n�G8i���&�[?�|����A��;�S��?Ұ<�ghPƯ�@߮��.��V���RVe��*~4H��9h� ���>���S�4��$��|�ӑ�4=�y�ܯ�+����{2� ��+[�ei�5@H0Ug�7��3���0��L�#K㇮܋?'嫄�M����҄�3_��|$�j��O��f�W�|q�s�� 8*_s�U�U�'��O:&H_�>�;��>Uo�J{�Ӣ�JUnRNT[	ݑ{X9��*p����i� 1}{�
endstream
endobj
3 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 4 0 R
/C2_0 13 0 R
/C2_1 21 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents [29 0 R 30 0 R 31 0 R 32 0 R 33 0 R 34 0 R 35 0 R 36 0 R]
/Parent 2 0 R
>>
endobj
37 0 obj
<<
/Title (1ec8b7e24be6c30b4bdaf70cc209ff749bbf40476b630bec24ca6359b02604cc.pdf)
/Count 2
/First 38 0 R
/Last 38 0 R
/Parent 43 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [3 0 R]
/Count 1
>>
endobj
43 0 obj
<<
/Count 3
/First 37 0 R
/Last 37 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/Outlines 43 0 R
>>
endobj
42 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227165622Z)
>>
endobj
8 0 obj
<<
/Type /ObjStm
/N 21
/First 157
/Filter /FlateDecode
/Length 2675
>>
stream
x��Z�nG}�W�c�@`�/@`�����f#g�����:dQ�h`��{N�5�Вd���k�}��[w�k�I�dB1����R2u��8���M��WQ{�up�Smt�{S�E�������g�ua�w���i�e���oФ�\M��y��}�X�����zs��|����r��}~�X������]6�<y��u�7����.�����������;>����_=;]���x\]�\o>��39����Z���l���7&��^�>��ǜ��f�W�Fy�??_}�\`?l.7�K����Q���b�s:�����6�7�_����j{4?�^>]������z�{��Y������Зou��bm�v��ͻ'�.����t���O0�|��
��97s���m1濺]�Pz�<]ݬ���Rȭ�7��忷��������I >���_w�tf.�`]��[sf�Y����/� �R�VP��Q��	1��&U��T�w�!q}�/�퉔���:�m
&7�w��L�N&A��o����	x�%���hq�'�u2�K4�����`Zq�*���^֬u¸���oų�?��<�d<���@_��c��<�[�n�sC��'�*`���	c�/XW�	k�6A�#�/���Aj�%���ǱMϯR�]n�L���
^��	\'�5��{ϵan<��� h�>[�86+�!�F�-�B��ሰ��LŦ�9�0�=�%29:��N7_`�J�><���2�}������|�ʻb��$�S�@���1(0",��tC���B2��a����@!��!�	I¼L�w�e
�{Ç����{�#O�Px�-�.�R�����E�s�iJ��@-������ �bZ(\�-?8[�Wg�p?�B��d�Q��)���\�餺v��m���|��V�R;�
$=�ZP�p�Rز��5ظ�V��>��6,iKk�Tۡ��q��LA�x����UFݏ'm����L�߭�T�{����t
P���@Hj}`IS�Pc?bUiX�H�Xk�J;K(Ϝ�.k�A�����&&���T�c�,D�����ǂ�����`�;{��A:A���?�$V $�Y/ sL�k ���bR����#.g��sp$��=�����:�U�PAS�wδ���,��Ј��lC��T���:��J�&2�����!�j�
�t7��7��ч���q����V���$MM��R�k�_Y\#�h꣮K,�v�������d�S���1q��1�Cw��
���8Aj�{���aO3b��:WG���˟��G�6D)"��cEA��ET{w]q�D;�ЃQ�-�F`}6FeC�o瀉܍�W|E�$�i ���级3�~}���ȧE�3���A)�}�w��`rn������G�We��m�sg�4}���G�փѯ�R�Mִ �;����Z��u��H�E��Xh�X��D���֥��l;�&��%�6½�>���Z6shؗm�}�t�9�EL���Zl��7��/a��nm���g聘���0��������Co�+�Ɠ�R�)('��^`�
<�L��-E��\a��>�{W+��OSa� J!��6	�1>�����p1ȥ;�S�,� iP�>��$��$�j�Y��R�8���U�}^�dQN �1���j���w2�G!sN�cC?��NU�5΁k?�����3�7�/����ϸs<�B����E�Py�h�P'R��-u�t��JCI���Sj<���H��:#�󄞻+�牪�� ��*�&%��ajJ�_r�@�{�z�μ�*�� ��5�Z	d�2��:k��g�\�M'QȄ�4/784�aHF��y��)���z-�*�!��#���\鎖؂��� �}�&9ۺ�#V��2 d���2��$��50�ޟQ�9�&�8b"*�&�����~�{}�gz�at�3y�������8❾�3Rzg��Ƒ/y;�P�J�!�0=×"�>�<%��`��� }e�~��O����}�o��w��ܩC�'�:��>u���R�|���Y�;Ed�y	ޫp�~'��|e�T�|S�K��煺���\*��sf��23U��΂iV���rǖ7&i��o��\�ɓ���W����r�Aõ�(H�A&��3�$��	�	omI4_� g��\�*�X��"��R��J�*�P��/�t<������P�E��"���b*O��"Tc!�kg�jt� E(^�(UL�Q�$��b"J(^\�(��t�(E(^�)ŘF)~x��)J��C��"#6�hB�Ҍ8�?N
�,�T�"�!)�
ͬR�E()B�BL)ƚJ�ح�J1� �:^�ՔRR�b�Tb*��+P�*�P�E����N�X@�5�K�~���Ձ����I�ܽ�����K}��0m�A�l_�z����V���}_�����P��t�˷Yy��EOFy���&��Ц�Z���TB܏�N���?ܰx��˔�U��2M��^IfE��_��Q��~$R�U�C��q,R>͊��)�����w�����m��,_l�l�	s&��ϛ�K�|��6Oh�u����������G��O�kr8�n�]�Ц����������w�6{�<�C�Y�i>��
endstream
endobj
44 0 obj
<<
/Size 45
/Root 1 0 R
/Info 42 0 R
/ID [<5217C64AF857029729064CF134102380> <216548CBC6346EF6CDBCF0B460D21CEA>]
/Type /XRef
/W [1 2 2]
/Filter /FlateDecode
/Index [0 45]
/Length 149
>>
stream
x�%�=
�P�����h�Q�#	��N,���&��`/��B�g��x�8�k>�va4��0_�����-Z"�o
38F�Iz��舮�-s�HDj�M�C������\8;U<z��eF�wrۓǔ<=y-H��6�ND!�bd��3sR��?���
endstream
endobj
startxref
50921
%%EOF
