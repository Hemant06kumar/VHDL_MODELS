%PDF-1.7
%����
12 0 obj
<<
/Filter /FlateDecode
/Length 20
>>
stream
H�j````b>�	  U"
endstream
endobj
13 0 obj
<<
/Filter /FlateDecode
/Length 1203
/Subtype /CIDFontType0C
>>
stream
H�|�{LSW�若�JS��5��qY�X��`�8u"�a��1�Wm/�(�p�R+Hu}���vT(>�<���XШè���8���l�͙�h�q������d��ߜ�����w�/'E��E_*���[���|���Yxn�j���j�`$aJ����(�)!|%L�(�V��f��D��t8K����j"�F^�*4u�����L��n���qU.�b.�3����tI3c� �c�FL�ҙZ�6�b���y1z���V�����Uo���f�֭L�����k����Xlk���<c�f��ϳ&��Ll����pR�_X�?�����b�E"�]\�1�i���Ū9���[X[��\}���e�[��抍�� ��!�PD��D�QJ,D~@�詸Yq-qc�����huΈf</��U����!�-Bh�C��9B��&%1$�I;ER��x�;�A� w$	$�6��50^'��,۝�j�YL�)��m��:�h@�o��O}�"t(�*����Lrp*z����(n�ִ��^G���8�qH3�Z�p�]oK S39{���z)���5X���a�R]���=>!�$���W�7���Ӏ~:z���@=�K{��@�l���l��[�HmE�H�V�K輒��s;$]�~r�$�q_�_ ���#4�D�v:��{��t��c��g�-M�fo�>�����J�Jv��4x�0�[�֦��"�T���҉�áχ�˃��0���6�լ������\k&W.	 �����'j˻i��͊N��!th��I�3[k$�/�Rh����=Ф<�l���ͻ�UR\�~3�y�~�F��z$��<8~��	�±Ғz���>.,jГ��;��iR}�1
�KMΤ'�`�8>;fD����c��\x�Z�vq~���s�)'���u�ҏ�v���P`�F0b:�����Q� �S�1�Ƣ�Ç� �woȥ���\���GUc�~�QHE���2�ńVH~G�d�q �1�:^�2��]��3��!�����EA���r�V7F��'���΍_:�;�G ���lt��(�7��n]�l^_�Xl�b9!��+��]��Qr�����/�|ᆶ��p��C�m�ZJ7��TRj��
i����gIu��nk;H���lU{`Tg�)������	K�<�  �8*�
endstream
endobj
14 0 obj
<<
/Filter /FlateDecode
/Length 262
>>
stream
H�\��j� ��>�w��l��a�6�C�д`t�
��1��}��-t@��|��7��>�Zy��Έ=JK��Y�@�qT��s�J���-&n	�n�=N��k��9{���&M�GBߜD����{w�-�����C���!<���+�h��Z�ʯ���S|�!�|N�#q�\��zDRg��M(FP��kr����nS�UPgYQ���"RuIT&*%e�+�Dϑ�,Q����	���Y���T,΅�q�1�Ki|�����+� {�
endstream
endobj
19 0 obj
<<
/Filter /FlateDecode
/Length 23171
/Length1 50404
/Type /Stream
>>
stream
x��\UU�7�.{�s
^���n��������"��������4o9i�?3�1�i��Լ��SZZM���dC�Sf��>��Z�8�]f�������#���k��ֳ��zֳ�A6���  �8SR�FT�r�*!'N��퐤���T��(�{����x�u���>$st�e�%��5���q+��#��D�1�%9剖��bB����U���MvB:%���O-������{j�2Ȣx�ۧ�*���l"�xr�(���3���(<�S�sC����%U3Si�q�zZqYnN�G��2�A����,�n������4�$���O&$�S��]^VY�Z@�c~�x^^�_>ൣ���N�����X30i��I~�'af"~�>�����z�6�ǭ�P�`��Do��q�+P=,)y�(�ŧ�%\�3� u,�4��t5Q��S݈�P���%, l���Ɣ�����ȿ�:���
��H<q�\Z�H7�J��	������<)t_ea
���I{ҟ9�.:�� �tͣ�IYD��d)j�P_N�y�2]C�%\#mH$�/G��D�_JN��w��V��#������f�&)��������B��9���#H-�
*�A�0YJ�����86O�������0?�ǳ��/$-��A��Kf���w�n�%��FO�˩��p-���tN���R���7D��!��]�R�熥RdC��P�
AeQCY�V�t�('oS
�1')�i_��r����S8;�X\סQ�Y�!�qȺ��%�dl��:�u��xc��m<E��]?�R�Ͱ��ǁ�W�
��@2�A�d����dz�"mI��G������R#N����\%��I�7�c!��0���C�̀ր���gq=F�2N���K�}�o���+!4�5^۠!A�l�[�P�1c~Ϙ�n�t[�3n)-������\�GZtV�Г�!�{[E�ѭdF��3��bHV�E�ꋻ �� �t0���k�>:J��#{1z4>���w>F^�l�nEL)L�K�j̚Lvo �i�~+@�;�L�EB�`���� �~O�p5`9�y������I�lm�5�Qp#�3YL�$���0�I� ��n�Kc�3ZK�\�� &��.��[:� ��C��F�����l���x�1Q oӕ�� T��݈b� �6�f�n8Cޢ1������9�fz�V��ћt
hMB�:�/ǭ�i�������+)�'���!f�-{,G|"��
sB�/��Pi�D��7���ˮ0�W���z���G��w�O�G�?��1F��j�gJ��Uc�F=?��=Q[����E�A[-IB��lC�(�'���g{��QK��u����p���X�b���)�B&�G���*(��m�Ӹ[��Ѹ.7"��0�u��K\ߐp�J�R�R����'[�\
hx�{J!I�t�p_���ǝ�q$+f.9O)|n�KH����-�:.���s��A��J(�E�t�S���?���O�IVP� �㲗���h�%�~�IhTĆ02��TE<��L�d�,�o�N�{�Jn�B_kc��>[��nz˛E�咧F?	����#~f����d��|�wk�G�dA�p��2-�Aa�|�z\��Ű~O�����M>����C�/�T�`;�'�z���"/����R�P���2�#v�S^Fl(D�ߒ�:�;��ԅݻ�>��w���Cާ�(�/�4�fG�%ٝ�|E�r�t 8\X�*"��ֵv0���aH�14�u���X���ո�x9��C�m��ٟ���^`̚-��/g#���<�M���5�RLf!�z��J��IXq.#e. ���<</���J����q�mݫ$� ĺ�$�u���B�h��*f�J�Ǝ�W^�v_E�"�o���W���=����3��Ԧ�k�������4�>	�{v��=��K�ԑ�i_@ ��U&"�&�6t  Qϟ2�@.�-���� ����"�x��F��t<q�-�E�O#�: �l+�e#������C�l0��!��>�Q��6H�Og��u"��Gω����Zم�x�*O��zgV��ǓQyJ ��T��}�k�w��R�mICi��1�,F6%�ݲ�T6u���?<��̄o��E�4ͳ�~\(���8=y��x�&"��.bn�Oy#�3JJ3@F��Ů6.���*�k��5�5�~y�r�\�!v�k�kD}<`{�j=W������{ډ��&�n��.��{�=^��R�7ݧ�e�RM@���zps>1�@�yQ���o�K�{��/����{�]/�e�Y~��M��#bE��P��������x�p't�����W��~�q��	t֠�� q\�G1����0�����d2����p��Gq��Y����vv{P���賛�$���>�������a�}�U���uyRJ����]��m%�H@�q����dD��D=г�y$�"b�@T��M��J��(�m��1ؽ��{Ë	v�IX��W���,�0�?gq2�ŽX;6�ɱ���$Ҷ����q��g�������i���{qh����Fo\���U���PK��+�Snhx��L���k�r���9U�[�Q�9Q���&Y x؍o�s�*�o�A���p {
�<�ҷ�a��3�!�p64<ֳ���mRh�<��c�0���F�nvw+,x�#o�Qnh>��[D/##�v�p�@Ns����[��܏���kEI|DA�����A��lh��(�"�(D�\���sW6%�_#�Y<uaQOk���&w���U+�	5î���y����D�bM
�e[
r���2��F��B�u���Q�ğف̆B�qY�\���S��z_Y����xn����<����Ç����u&�����[���ǅ��J�������x�URĝ�ɧv�  ��L�y[����Tߖ�&�D��2g4y>�����O��� �~�p�t8"h;���"J7����G#?3#wΕ�����yG���ؑ��A!'�Y�z9](Z��J�h#w#����Lau���!�]0bU�j������C,��Z���j��n֒�As:NW������$�V`o�F���?B��w�g8N�pJ�L�;2�h��0��ݐX��B'�j��Ԃ�DE��@	G��8=��^X�w�A�mwĿ�(w�eF,�In!2�x��{�S8���u��Zm�F�$6%�n�h�6}:�y��F-r��<�Qo	��'ZCp��V�����V,���п ������pZr!JD#�%��Ur��Rd�I�-�_��4 '�LR%Kw��L�>�L4Y����>t$�8G��]�b��?�8$FU��]�{�s:J��'�մ�L����ȵY��4h5v�j�FA��%�1�#�#0�n㩫`�1�?M���g��K*>?ތ�G�'��$���E�Xg�cJ�? ���c	S���B����/�{.�u"�n-W�������y_�I�g�8�N�X]e����uш8�H�zP��$Qx��*�;�X�1(�O��%��>�����C�Ok��c��-���_����AOr�:���Wdl�M���Z�k�^�\�ȫ��������0��ë�B!�G�:W<�t}��4��If����N�ŷ&��7%����d��0KF�6��IFi69�x7��~�3� 7���|��� �$���i��$d0֡���c���Wd?E|�%spBN߄ѵh������I1��1�p��hD�2+1�L���,��G�r����� 3�@��C�ч�\�/~�9>��[����%>�;��|�C�k.�5����<aD|��7�Ǣ܃�e0J
JG��"��Dg�8�F�Mħ�F�e���Lr�D���'���2�!Nɂ]��I����a��R��HO�ר���N���-���]�Ț�&!o vɖ������E��8�;x~:b?댈��#4��Ё��.���L!y�/��P�ð���'"��D�����au������������;<�E��*�t�ӱ�E��퍿7�yj\��Q�n��s/��g�������Q��U����Jd�g?���Q�Ge;kh��$7���Ih��FUܡ��I�u�����:s���",s����O����_MhK��	s��D��DG������˺Cb?�	�W�}��c��I}�pjG������*�Yd/3�4NM���>��+���&[h�8��:����t���o���7����P��G��ߏS�����+�_�~?��\�ȿ�6F��&�6��K�Wu��8~%���ׂ�Z��ָ�ǻ��__�S�^�/��t��/ۨ���m��t~����??�?�4D��&�4�����t��A�:� ������� ��:o�M}/��;��3�_�������~˪����������e��m�-�_t~v}y��������\~J���U���䣞��q���+:?
zG�;?��A���_>t���A��|���H����P�r0���K�xͪ�E���e�M�g�zA������}�� ��������:߭���]:n���\��˟��>ۙ��������?s����w:ߦ�gt�uK��5�oyڡn	�O;�o�|�Ο�$O�|�߸!Zݨ��|=�_���{�N�O·�<ȟ���]������W���	�?����Ց|��*�?i�+m|V���P��H�̟/���/������Gu�ȟ?��:�?Q}8�/����|�Cs�y:h.����_>[�3t>]��Uv�ڏW�P��Re�UG�� ^�T��7:/�yYi�Z����tVK3yIg^����4���|�A^��|���<wJ����)ġN	�9:���I:�x�M������N����qxtv ��1:�&Dǳt�����;�����@�����:B�i���|Xj�:�/O������P��ݐ<�����<9�'�!�/����kX|�EIL�S�yb#�K��U�xB=���Av5ޗ�����d����|P���S����`��|������?�?����Z�7���y��j���{ŶV{�=q��8t��y<�њǶ�1���hKK5� ��B�Ȼ�01m��_�j����n]#�n:]#y6@���:��~<�e���;��������:o�쮶�˝�y�p��Cu�N�m�۶:o��	�u��`���V)�ePw�e"
t�A�y���@��< �t����38���Н��]���~��|}��������|���{A�[�]�V_Ŧs+$���Ғ�ܤs�5����C8~�Cw����88��y�V�n����n�g��#�Y�(���Ѳ��C�����*�����Rz ��x!��Z�k���Ā�Ri��U����U�駱"o�<�j��9�ҷI{�	�-m�������y6N%d;��s0g��pe���[f8�/�!�Iꂳ���#��$��v��8Ϝ?:�_9��,u���f�wVa��D�S�l�:�L�Ⱥ�����)d�zQ� ��E�*��N��M�B�m=D{�t�6�d�	�7��H�Pf��d#|2N�o��@��AVit�2Y�!��L���eМ�o྽�!1!/�5]M���w�^e`�A��oB�3�UR� <����
�ad'h��2����9�J�.@wu%_�R�'�)�����:�YƓH_��N�B��71�%�*��"�/��)��v��&vH�Qǀ��Ԭ.�Y-�ą��q��Bml�������*����������{��
M&�f�]����!�ӥ
Yb&
��
J����R�	|ޞ�{ԋ���(��]���Z�Y!,�O�L���1��`�/H�����*u��TcA��":�޽���E.ں~���Z�%��/����
=��'�D-�N �N�&A�Dmf��@��6��nϖA���'�w/F'H�[A]��~�>��+����⬳�S����Iz|���FWM
S�������V�.�l�r�揬��?�f	����QZ��h%�&ZN���Rj����N�i_տ���M�D��{+���i���?UIG)�;>�u}1������r_���ů����Ox	[{��'[�B��pBZ3��jO���p;�^���!B�~���v�/�#�A/�����D����P� ���j�o����>Ծ>x]��A�m���M�_h��P(<�q�^���+�����B�Qb�-�c���Xcl�� :�⃔A� m�i�y�e�u�m$IG��֑�Id��&Y'ٶ�-t�·([�-��������y�<{�?�<�>�=oz����y��#�=�#���v�t�|�r�zĖ�S̸�ⓔI�$m�i�y�EL�S�:�O什��k�E�wl��=�������~1�O�Q#���h���+[���~��?�y���wԨ�����f��~Z?������Kc��3����L��>D���X�X�DI�z����|��֫KLd����rX����F��&0��;�����/���>u�v)�i5�n^�E$����%��w!m#UMi�[���45�������u
Yψ�ʨ5�U��wh��\G���wOx�l,�w&�������*n\x$��݇������1"\3�����S�3�/��lO]�A�;/e���ʧ�������wq׮]'i�=�׏��X��=�.�<�hU���m����v&C�o��A��>뵰��m�G��6=ץe�CB;:ByxX�%���j��⫅{
�~�q�/�*�b�ޡ`�x�F{�&Ls���?����ԂW��طoæM�7?��Å�^N}��KyX�מ|�;���k�ʇ7�]R9�s�N���]�M�O+e�#CtJ��>܇p�H�ʹ^�|��ڭ$Ԭh~����:(���/�Z@C��i(���pm�{���}o��ޅ�����^;]�XmW��������4���*�;�nG�WL�Z�7�/w<�އ�'K|6�v��P�*�ZÉ#,T��{=_r�K?Z���B+$(�4Q��כ�Z��nc�����f�L�p ��?|��M��]��?��׵�U��/q=�nۺ/2��ę`��E��B�[��;��W��=��o�α12<�t�	7imi��Hn�.�����s�ÞA�T,?���N,E�>�%ׂ[��O=6�諱�J����Gzݷ4�[��`���.Y��p ����������V�N���t6]V_|`���Þ�r�,�=�B���F2�x��*�*4�UNN�L����tb��z�(�¡KL�~9�]����\�[�8��������t{#Hl'�;i�C��@���\l��C�Р�~�Р6�<ԯ}X,�V+�&��qwq���RAd4��;���k�ZZx:���p�'-Y�~f��ߞ;����m��K�tז�g͞?oά����e�6�_�tCV���;~߼ڷ?��̥/No=M��|衙��/0�dJ�2u wŇ������w�,�?�X��o�.|cd�ӰpK��c�0�ZXڳ����V��y��� _aw$=����Yւ5k`�ş	k�����c�|���#u-[�1e�R����!yP�Q��L/��a"ב���I�:m�}�6�[٦���B�rkA�y��7к:��~^�/�Q�X�ƾ�XHd|�6���l�v[�B�QS;͊�pVZAA-�G��������r}�+Ǽ�/���k�y�{�d�2K��k�*�����`��tV:	����F-R���2�n����=E?��n�A�	�d���,��-�]٪��ĬRC�qy�X�(8/2?~��Y�.r?��HU��?�4�Y!�������MC�����'��'�H�k
>�>B��[����k����ɾϱ޲�ol�"�Nzh���|���	pc��r��/����m���~����o1lט�'N��~.�w�.t-��tc�.o����/�������.�����6#�����,!��4�g1�8{S�#6 �ԉ\U.p���>����#�[Hn�P�q�9�"������w��w�H���?�8C������?)Ru�S����5�%��&�z���?Z�j�aB��i�cO�I��"�I>�>�=V_����17eW�����d���t�o᦭����{Y�d#.��	,����š���Jzc@o��ɢ�(3�sf��Z��V����6�b挪VMSb���1�&���
������ͳ���Rr|�l������9�ґv��],}p,�c�g��3�iY����T�#� �a�~������af7nvS;�}�[��+�[_���o�[X����A��6�8{-.�w�d�~b�'�C�i�U�Koڸx��M�������uH�/�T�Z�RQ�ѿ�!4U���GN��.����ҿ����� ���z��%�25Χ�?	���fq�K�w���#ۋ�D�q骯W�v�J=��p�2����gԘ�7�.Z�f�|�y�N#���s�@�7-���l�V-�+\�T��)$�+A�-H��տ�E�V�O��rkH���#�j�mg��`ʿ�D�����9_��G�ժE���Wɶ� ��^���_�������t�u�=S��[���X�C/�����~�z���d��<�肥� �rX��W�["�6�9�d���Ōd�$�X�%�H�Tq��Fl4�[�ͬ2�i�lf��T�ܥŐ���X`��.5�g+/i��~���ڗ	g��*�`��̻�mٶ�l�:�f�e���́���=�T��#m��h6Μm�g��!����_��1E�H���@?����^�>���Y�Xw�-���[�5X�J�9'��6��LC	劌�"����h$8\��z��%��ݝ�N9��`�ߟIB=�9�>1"qW�����e����"�9"&����Vi�����`ӊ��˝Gڭ�p8`c�VB|��=ɩhA�tE�G�g��cN\�Vw͝���Ip���o�m��l�[�V�V۶�[[m������4�����?����;"Q���!ޝ��D������fo�C_z�?�������>�f������������My~�����/ؑ7�m��{tV�^5�:edĭ1d}�fk���-��ol��~�A��y*�	�kZ�v�-.�8t���/R,OV~��A�q�c'��=��%�]���EK꿈z���W�_��]S�b�y���>|�����q��?��c3W��p(9~"���ھ�稃,9�rw��b��h)�ag�~�Я�<�6�G�J��f�u�4�*�nJO]s��=yCB�n�h?��5ꕄ��{��z�>���ЋJ[��\a��{�>�[)DcC�lC�^�ɛ�EdF�vF�lI��L~_MM�Ƽ�/}&��dѢ��-Z�ϳ���]�9�ޅl������y��?x��O6�~��;����4�Rk��j+|�+!+Z��؎��KK���p�y;��o��pFǵ+�Eqvh��O�Gs0��p3%��#{�������O�W���Fy|ɢ�6�>��S������-�����������~�Q������v�~�� O�jǬ���XT���(�:�Zr�\�I �{�)�ގ�]���"kW:��A��j��s�7�;5wU]?�*�f���s��J�{���bm�����hiY�r�Ǌ�;��X�N!D���ł=��}'���xEh���d�ǿ���q[����[�`�c���[\s��i;2�l�䒨%'���D����w�}�Ϳ��T�׵m�?:j�^�܉� j�f:`�}�9��_����`�/�Ү�?l
y�F�� z���(��@d.�����2-�ABi�Ҵ�,X^S�cg��c�뇱��{��������s?zۇ��0�g����~b?a}���~��٨����V�/���@�Cw�.����H�#(��Ғ�RZ�F�jj��u1�V�D6���k+�ja��#2­��'�~�c�li�h�Y#���e,��]�:�~���������W�	]��C�/��^�%�3�=��.�Sp��E1�vm4S�}��ns,�a"�~�Z������#Z'G8��k���?k|�K���h�que�&?�8��5�A��Z��X%V��bM��XK�5�6��V���j=�͠���
���+����|�|�|�|�|۪��Z�
^����6�ڮj�*4��/�d��e�F�ɇl{xѰ�e;{���kg�a���}�}|~eh�y���l�7�s�V?�-�Z.�����4�t��w���w.��w�~�w��;���b�P��d>�� +�b_��%�{�e j�'�N�����W�X�z���?\��������߹���y����9�2o��4IU����>F�¼"6��o���n����v��Cd��ڵ���sd������>6㥗Dx��Wg
6ҫ��=l���ӚuU�X�U�klY�����ۘ��J΃6���}����6�C�������4��<y��ipA���xѢ�K-Z�Zwߘ��Wg�����&x�Q�,s�]�%06sտ���ɧ�BO�d$�c�q�����3�hB��'�yL\8+�=6>�A���$N��%8�;b��I<��EF�Q�Q��Sc{m��V�»f����Y�4�������o+�?�1/���.�_4�ӉT���ؙ��UX���L�V�a���B����0%�,�G���AG�W�++"�o���jkc"#�h��&-0<���/�P�����"h%S-���t��I���0�A���y^�|F��2rk��9^�te�[���M=�5�����[�x��};��/DGߛ9|X�o��sw��8ܻw��=�oؚy�<�^ʺ�7�Oc-���U�~|?�����f�����t��6����R�M�?+��������]bT�֏������5;^g�W�{ܹSeb����J�����  ��a�8��o��𾆴����^��K=����t� b��Y?nۙ���a�<�X�L&ɏ�Vƹ�g�ޑ�k�8S�'$TURI�I~&"��A�N�`�k"��YQTɘ�@#��d�rD��{L���V�w����N��m8�[-Vq:�Y��<i�L8��I��$���k+bO�����F���v��b6~c�f"1g���9��r$¹��.^��6�b#a�k��*!j[Kkk[��#�i�uT�h]L�({�G��7�4�'�S-)�a�1�l�X�8{+�J�:͒o��f�3�Z*l���!,���h�5�ڍuS�a���C���X�Zh����Y�<e���u�5z��ن�4�F#����m���7��i�^(pK�?̗����o2�].�.m���j+ͤ)��bU���Vj���V+�ڵ��n�&�*f؜�k,լ%۱^�N���~�!�$5j�������Y&�D��5�:@�e�Oc5CF��I��2Q/�5�����F/;K��N�����k�+� 6���'Y��,��dk|�O+_�:6f������
 �V~".�_�V��>��>�ײ�t���X��Έ� s@�orq4�{�+�����*�?21�Pz|k�1�����{�OGߎ~��S�S��X�'�C��K�/l�
I�wF��^6amɽ��#��4:�8-�>�����i�	%�n-/6d��d���� dz�$���LVǅK�ߪygw^��'��{^��> �#�i-=�k��%��oUW(�yJy�z�a�B,�B��D��H�O���d"�~�t3��Z]$���_| ��}'�z�">�y553^�����5�O�<p�8������:���Hb|���}�����1;U�,&)�̈́��/��'��dKr����ȑ`��l��F�C	N'��/���U瀙�^�tl��^P���� ��ր���Ma����.����lV+_��j��� ��Ӻ6�e�3&0�j0?����-NK���u�u����k�ٶ}�+�~���g|�}f������_�߲;���;p���w�܁;p���w�܁;p����灃9R����'BZR߆�m3�x�Z%�uFR��Wl���J��]׈/�箋���]��v�iw�ǲ�����^h�*����8m�:#f�`w�{�+^u�ۆ��ik�u��$�6�]���g�u��wݗڞ\V>��hja��sng\llO�Y�Ģ�ʪ����(gjin�3��ؙ!zU:3�+�+���E[��匩v��Nͯt�T�;�J���S��r�ye%9E��>�9���e�e�ee�ɯ�,*+u�E��k<��SwRLT��������}zuteYuEn~AY��������E����ό./,�I+��/��O��7B�I��+��S��ft�v�
ޣ�����9�iPnИ����X���n��f.�Ϊ��������eͩX���+J�*�bѻ0�"sM��)��ϋrT@x���^���̙S:�YS`@ٔ*\T:��iѳ�0�m���ܲ�rt�
A��д�s�TIx�s�TV���`>h0��$��*�J�SPTw� gfYA��<���"���,�:7_��+�`ES���%MD�J���y��EU�e�U`���=��_a�d�+�_��,ɗRK�VFy�%�)�pV���]V��7�Z0��B�Un�ɉf���:@������ˁye�ʲ(ge��i��U���q1\R�[V�W$�`�f�QΔ���RË$NPZV3T��*�`<sV�@�)�n��8yN9�J�Β���ۊ�U�_������>-ə%藔�	G�)����9yyRrCub}�T����
9Q^~e��R����Y兕b��М\�#<�T6���<Ca9�^�q����H,��r5qu�T�/�%��J�P���g�����f�U�U:��b�����.�n�T��N��IP����ˊ˟Y�U��)/�˙R�/�r3��T9s*A1���^0]���9�"�ƕpC�leY�X��t�P9�bA�^<�srș
��K��ǯw�&S!h�������dg���,g�Ȕ��	���L稌�cR�����	���r�M�:rt�=2ҳ�9G�8��9���'E9��Ge$gf:Gf8SG�JKMF[j���I��C���>2˙�:"5D�FʡnR�ə�؈��Cq������5.ʙ���.h��h�sTBFV���i	�Q�3F��L�$�MOMO��,�#�!9j\FꐡYQ���(gVFBR򈄌�Q�Ñ9�)�D�K�p&��3�&��9S�2�2�F��B;C�G�:�����:2ݙ�QӒ� �ഄ�QΤ�	C�3'���4�C���������<8UT��Ԍ��Y�'tM�Iv�L�L�w4��324YN�o��L��q���Y��M�L�r&d�f
R2F�]aO�2��>�����
��[���h��I�	i �)ظ�/�+yfn~y��m��6£�F���^k��R,\�MV��XYr�1"\��[r�;�����nd�߼�����"�`}��`2��R�tl�%e�}�2��aTC/�˜b�l`���l��E2���
�ęS�֊��½U5�@�Ҝ����r�TE��gE�o���$'E���JܢK��V���*�TI<�#W�vZ�`$��d� Ed*)$U�I:�\��8���p�D��Bb]���$���(���R􏖯�)8IF�Jy��k>�L�CO+IBm(�!�葋�9�2U�t�.�;A��}��n�91����g��dJ*���*EID)#๘���$�8pѓ�m2�3�3�)��jHT�^HX��?W���?��ѯ�
��1�BJ�Cf��Pb�$b�L<-�r��Ii�%?�$�kn�n<6��&�Y�����n��\f�"-��F�������sj�<��cV�'��[����[�/�\�֢S>ϑV-�Z} me��_�EH6J�+��=֠](���*g)���'�ȧ��6|/J�U&9,���ݫA�¨�m�"��,�nM{hVI.����B$�!�n�
���{q��
��pi����K����n�g�`.��DR��O<�)@���ǝxl�AD�ւ��b�F���r�2�R-�l�&OJP%}m
�Vɧ�9~z�(�Z�gՒ����
e��rk�D�yK�_��+n�����#�%Ҟ[7��J���	9�䌑Q�))���]��jS�����ܖ7xtU3�k�h��Gɯ���
d�-uK��5c��b�(y��������ۏ��Q�c�\9w����� �:�ܣr@�LF�FxǢF�	��R�^�M�z�J�mc��8��9�m�)q��k�6�H��3�,�;��m�y���-�̒��( hG7��ύ:����\}Er-{"������S��</�{{�g�����9�#Q��Tث�KS�+��.\�0�'��H�1|�3Gs�T��L�1.����Hݎ����|��r;��v/��~&�W�#P�䯤	]OKe�gz�M�]$���X`��*O��;� w���g���6c�5�g��u_��k�{=x,1O�n�1��U��ѻ`�b92��7����ϯ�B��Z��1_z�O��!��b�xZ��"�����Jx��k�RFOϞݸ�<+Jd�9H�{DS��ң �궘�/�J�6�?���X?-���r��J��<#I:��<#q�E�"�̐��+O��#��T�']��<\�Ʊ��#�hIˠ�,h�C�����n8�����,_w"f̔T��m��4\�����B�Ѹ�!Dd��|��%׎'x18�B{�M�J�3z8����~� _$�&i����zz�)nN��eAs08J�w�u4���/S�3A�lp�.eH�sC�dɁa	����e�d�,Ʌ�)��3JJ(�I��Ŭ�e���H��E��J�[�B�cfΔ��R�,�"a�������IaD����%H=��3$�gB�B�i=3��2X�K�Mp�$gJ�ɼ�$jM�s;���0Dʗ,5�&{gB�����b�c��u�[�M���H���`)��콘5��S	RwM�0V��Q
�	n<�Kg��Ow[wp��GJ/�U+c�ZL����3��"��7磽<�c��n���YS�z֑�߯�-��M-�$�)��af�6~��������󎱯���t����R��3�4�Z�L���Cdߒf�[��l�Y�g��v;��l��ٯ'�0b�q6��~�d�n䂕Y���5d&3���=�8����J9�!Y�{DsZF~�#�1[�m��s;T�b���Yf�z�;3�U������N��NU�d�,���
i�rb�����E>�[A<�F����4�z��	jH�<T�`��yn����9�����C��ӷ}C#f"�@d���e��=�p��P��mDmۄ�S�Է�ߡ���D�9��߳�Q�����G���Q�_a���{�S�꧕9�**�	W�(o�~N9��y�-��V>E�3�g�ʷ�0�%�����_$�^�.b��G�k%{��%��e��99SHlbr�Ԋ�Ȩ�2'�P�SU�î"5ᒿaԘԐ��̌D�0�Q���L��E/bN��$��K�&�i��.>�'�2�g
,[(��P�8J�^%�<@TTMɓo �����P#&)��K^J,�%	%�[���ě:��jsd��3AC\���t�qoyи�>mh1��6�����'T�H�=�k[�D��٥(+��$F+�J�@��|�Pr֑����-x��k
X�T��IyXY�+W�)��3���?����W�5�)���(�I � i������3�O!=�≧%օ��nׇ?�g�k	��r=�в��Rg}�,�d��������Ł���>J��)���J-yc�QS)�Ъ���O间�~KoP�)���%k��Yg�z�,���4����D�Ǧ�r6�=���|������v��l�a��	v��c����+v�]c79��� �Cyޕ��>| O�Cy:����ɼ��
>�?����j��o���N������U~������K�k~�_�u�/�+�J��Zq*�(%N�ܣ$)ÔQ�e�2E)TJ�*e6����ByB٠<�lWv){���!�rJyC����|�|��*�*7]UT��P[�m�p����R��j���f���D5O������Շ�%�c�Zu��Uݡ�V��5�a��zF=���~�~�~�^Q��75�i�]Ђ�P���U���h�Dm���ei�i���X��fji�h˴��:m��M۩��^�hG�W���[�{���%�k�v]�31���k
4�69MMQ�8S?�=�$�0�(���:[Z<���������	Ѕ�
?cU�l�u�g�o՟X�"�����+D��O%��Ҁ���;�;uD]��*.v���Ւ�Im�l�J�'��\y��6����:��,^A`9���W�W��W{���^�w�T�͖x��-���B�A���%V{�ē]��}tpΊ�w�H<����H��K�%[�8[��8Q�L��aI9M�񮧀�sm�uђ*�Xْ%�ѳ���e���[虮u�_�O�L?u�^"��>E�*����n]D�l��d�P���KD�l���~�Ϣ�Fj��_(��d������1$�zU�F�[z�6�yLkd�!q��� m1R�&4&�Q������J�/�YZ_z�^����8I_!98Jh�#�z��U��#R6����ʖ,W0�_݀�r�����T�1��I���Mr�}[LՋ��������CRB�ٺC�3R�%:A�6�Enh7�L=P̥�7kO��^���U����7���Q���m���ր�����ڟpm���.����]ըOs-c���_�'(�l�k8Z�w�+���6��҂%h��Im��j<@�ܭ��0�$��I�|���X��r������t����o��������������� dV`��b���͔�̈9I��5��Kƙdi�!�[�LDF|���X$Y�e�^y��#�#=���HRf�l�F*�w��"3���d�=ž�̶�F��O�O'�O�.�O7�(���ӻs�7~6�٬	K�1�n�2�Ҭ�)���<E���t�Y�Oԏ���	�e�li�e,���ʌ�ae��y��-`��O�T��~�x#�xc�0b��si��݊���R���`zЄ,��x���J�ҷ�{�cz�~M��봎1ff�,��fN֑E�8֏�Ò�06��a�V�JY���G�
�����YeN'��!v�7��>��}�jٷ�ӹ­��[�<�w�Ѽ��y
O�<�O�y|/�����a��?���M|+��w�}���'�~���?���~��T��)v%@	VB�JW%V�T��J���ܧLV
�b�B�	/zDY��V�)��m�Ne��r@9����U�R�S>V.)_+W��J��T����U��Q�R��~�=j�:L��Q'�S�B�T�Rg���G����iu��Kݫ�W���S���}�S�K�V�V��ꚢY5��Rk��k��h��6@��R�4-C��&jy�4�\��=�=�-���j����m��O��k'�3�9��C�s�+�vM�i"&�$v����yf�ϩN�ֳJ���&w7V'"���A~����k����"�#E��s�؅��"sP�(�A56�_E�C�i<e�KA�:��.�H�v��zMD'%�N\mVo�������NHnE����WeV�E�٭�Oqe�d4X�~G��&	>�.�-�"/J�x�^$q��Y^x��$N�x��yY�����������8Uy^P�-Y�)��(�pU�����V�,��kB�Z��d�S�¬\jh�"����d��>�wH��-����E������$>���ʔR���]����Wa�GU�J.��_�&�I|S���,K����F��~�w^�B�H/�^g7��%�,v��(QE�+bi˅�D�b�KR�wi��(MP(��L��������Ke]P@����D)'d]��\��Ş�T�$�,=M�|Ax;��>Y��Po�:%b"�UVK�~.���T��8e��=ή얜�B�,PЇ��l�.r���~?e��������7����I���yA9m�\wvu��g�
���S|��s8��΂&9���K����Jd,Bo���\���%�����~Uh����GT!�NA��P��~ �}D���t�&�?�ha7�~w�B�b���'���d����Y�@�,�M�����ŪJ�
���biy2.����k��"J��8��D/	���<CXPAF�x5-_m�8>��e4��E���o��wAK�Ew0�T����3q���S5Iӈ�e
��m���Et�"2?w3N�9�d2\yFy�D�D�,� ��2�ɓ�L��g����H�=	��o�Ʉ��|:!��X�3��|�������k�ҕة��Pցue����P�β�}l2+`Ŭ��d�G�2���c��6���a/��٫�,{���>f����*����㟾<���NޑG�8ޏ�Ó�0>����^�Ky����G�
�������.�����1~���/�����K^˿�7��(�Uq(-��J��Y�Vz)�x%EIS2�le���LSʕ������1e��I٪�Pv+���rB9��S�Q>T>W�R�(ה�*Q5ծ��j��A�ƪ}ԁj�:TMW�����j�Z�V�3Շ�G�e�ju��Yݦ�T��/�ԣ��Y�-�=�c����zU���iL3k�Z��Zsj�(-N�ݣ%iôQ�m�6E+�J�*m�6_{T[�=�mОֶk����~�vL;���]���>վ�j�o��nRLV������n�l�6�20śRLi�S�i�)�4�Tn��,�a��c���M����ݦ}��a�	��9�;�M���2]1]3�4�f�����PssWs���y�9�<ԜnF4P����?	Lg��lY)���R��WO��k���>��Ю��&�܂��[�3���rΫ>ݛ����{���>�C�KY�6��ݧ�uL`�5�ѿ	o�����%�yl��6�'���4���L{y�|���[��⟝�[��%�R���[�n�����l�Os}�볽$�5�M����u��>oԃw�?ֆ����U0����qs�UW�7�������W���Dޫ�֕��b#J���s����_��?�W}n�/y��bD�p�Ϸ��	=7�Wf��z۱QR�o�]^��\o5�D����O��$�o���oϑ�S%Wc�xt�x#9���5y�,&��2�� �ȳ$��"5d,9@��r��$e��7��+� �/0�o��-��<I���zr�ԑ��E5��Zh�������5#��4��H;Ҟ�%ڇ>@^���ߒzz�~O\��@��Y۳�ٞ��?�]}pUG߽�{߻�~$H#Z)E�0���@i�1ELc�!Jhh�i)RDD���4b���i�4c�0�E�0� �#""RD������e��?��o�/����{�9�{��I^�!�Mm�au���������S��E�5�^��ҶH�UڠԱLJ��Y�/{�!��s�
�J������:�^^+7�-r��&���.y��_>(��˝r�|N�(_Q�JT1_�R�(ÕQ�Xe����(yJ�R��*�J��HY��`LY�X�4*��&e��]yK٭�U�U)G��)�r^�a�>�ؑ�HF$32,2"������X� Q���(GT"j"�#�"+��Yd5��ь؈،؆��A{��C��E#�!�F#�#g#�x����@��7��ng�Q��Fq�E[��7��-�����hs�
D����rD��фhA�"�툎��<�GDAGtF����xq�15���&���OES!� �#p�T�"& �9j�������! ptP�Nԥ�*jE]Ce����[����ս�{��zB=��Q�#���9�W'@6"2D~Ȅa0����8����4@=����g��5���JX��u�;�;0�I�P���p��I8��,u�;u���4]s�tm��o'��´�jN�&L��M���D�^O+D����jN���;m������wԝ�Vk�Z�Vu��δ�.�MC�i�7���޴ND����.���;u�c����tԞ���Qw:�NG��;}�>A��s�<=_/�K�y��Z_�/�W��5z��^ߠoҷ�������^�]��~T?�������K3�`�F��adÌF�1ΘhL1�Ӎ�ؘc��F���Xf�4V�:���hl6�;�����>�q�8f�4Ng��eS2S7]3�h6�4G�c���$s��k�0�s�YaV���s�Yg֛k�&��l5��v���e�1���#�q���2ϙ�+V؊Z��[��A�k�5�kM���+�ʷ��Rk�����YK��*k��h��6X��-�v�-k���z�:d�NX��3�y���>6ض�fgؙ�0{��e��'�S�i�t��.����v�]c/���+��v���n�7ڛ�m�{�����>`���'���Y��}ّ���Iw:��;���g�3ə��:3�B�ę�T8UN���Y��9��Z��iqZ�6���pv9{���A�s��t��s�E�v����nw�;��rǺ�l7�17��(B����.z�������.��.��������.z�������.z���������Q���S�3�b��CK�Ћ=�b��Ҽ/���q�Do�7͛�x���ܫ�j���2o���k��y��Fo����������y���1�w�;�]�.����������������H�?ޟ�O�s�~�_���+�*��_�/���z�����~���w���=�~���?�w�]�9��%5�M5S�����R��F���?��V�YQ��|��xl��D�)6� ��m�����ڞ�`;o������������s#��y5ɫ��rb�<8'#y�ޑ�G&��{+?�w{/�(?Y]����]m�^�Q�ߓ4�����Z�ak�z���뺒�AK��-1�|�ܓ4+�Fvգ�s�6�5�}W���M�+��D_빵��u�b�C�[)Oc O�gcm��<�Ǔɓi*(�c�lbpw����٬��a�6��ڹ���A���-��UA�ldI�' ��<��"0"G���S��60���H��+$	�����ډ�XOF�d�[��$��Gy��_�zBkH&�g����]	�����m&�=޼m�g,�m����J�	��(�y4�yg#Ω��	y
���w^Iy*�A����T���H�E�_A�"�l����$�s�O�<����3�xnlU��Mړ�� o'�N��.������gM�Ϧ��"+�s&���E|VB��8K��kR]x�I����%q���f����������n�C&��I׶o%��H|`���'�N�ӓ�9���m�M�bW�x �N��6ݚ(ORW����JݞrV�tGψ�~�3�L�Ø+�=y��?@��Eċ�W�$���ji��y������L�3��/붜 �L|2�~����ڬ@�]o�؃2�$�)b�M)��$M���ӛMyf/&^����vc�2�e��Np��^p�I��2�e��<wS9��4�3�Y��O1D2�3��a%`-��v�}���v�=l!��β���#v�?�^���O*�ğ4�����%�����%O��J㥉�D�$M��������S���ӡU�:�Bh��j�RRSR�ꔾ)w��S�My���lO��_�'˓��N��?������zyUn��&Z-������7���m��V��j�6���qޮ���O����k���WzM��2(:k�e�AYwӮ��W�"BE�U�S�3��K,&$�� �F�!2ا��t>�s>1G �whB��)��8&�r��*>���J���Ԁ;��^ �f�w	���ւ8�G+I���Zǰ���ӈ���z�O �Y��gzck�����K������mEX�g�J>'�H񷘄OX?
D�eK�rV��ы�Xkem��u��a��Av�g����"���<�M���|�Q|,���y�������y|���R����kx#_�7�M���w~O�M�Ů���{[N����?�	��K&�E.�qk�7LDJq�(֒3�!���b��TD.B�Y"J������W�X��b7`=��[���:��ykA�U^L��@Z|=�f�׷���>�a?��Iq���YBq��Y���(�3%g�P<e,�Ӿ�����M#A�f���M��x$����`Jq�Z@q�:��B(.tŅP\h��������#q%�o�Ģ�f.���Ϛ��6����16uNY�L�[VQV�f�`&+,�?��\�s��]Z�**E�*�����O����5�P*_m����)�_eiL���l����cM��K���X�]��+֧bG��ӱ�ãT?�����
]'��*���>���rE��8^gR��x�$���f"z�~�>�L��(>9����L%����X�$�#�C�
�iO#��D9�x١�~��U	�MyR\�$�h����~x ������"<
_��0�2x��'�k�4<�·�;�=x^���ex^�����?�?�Q���"�X�
��_����`(|Z����Ѐ+qFۗ�Wnӆi�p�"���v��#�%�2|f�|XO����M�6|������~?���u�?�?�?�U���T�� G��� ��!�k�0�}@�(\�Y.E?,��"b��Zl���X���?�4�vdC��(�"(�
��j��Ű��JX�� ��Ͱ�f��zN�TO��3�>���^�t�k���e�A�A;�v&���~g���z"W&ك�\؆g�-��m��s�̛tf+�y��|TJ:yEшxu�y�٨������w^�\	�ϐ6\��b�Cl{V}��������]C��q��?��o
endstream
endobj
22 0 obj
<<
/Filter /FlateDecode
/Length 457
>>
stream
H�\��n�0�_e.��k��%����V��8)Rc�C.��5>Vk	��}��4�n�s�Lū����8����x����=���~���;����]f{޹�H�5oa�2��=�������܉�ޛ}���4}ڳu3�T���c��K;�mϖ�h���a�o���s��m�TE�	c��ej;�[w��.�U�z�����+���}�>��Te\JUA=A=@5P+��c\�
/����PA�K(a���
6P00 B���00�@��(`�-T�7D���0T(+S�PVʼYR�͒:o����6��<��r@�Z �����!4���!4
IPk$>�a���)&��SL��z�G�ME#��~΃�H$��I1�dR��dd��Z$�B�B�7Ҭ����XFg����އ����8���~�)�qZ\��` a�c
endstream
endobj
27 0 obj
<<
/Filter /FlateDecode
/Length 14941
/Length1 35396
/Type /Stream
>>
stream
x��}xTյ��g�s&�B!�W	B��~���$$�2�LH �ę�����R�R�)E���H�q��Z��Ek���T��Zj)�3��^��d���~�~�e{�}�c��^{��3�3ƺ ��5mZ���3g�`�A(�==/�wbEc�ٸo�^R\�����)��z������N�y��[] ��˺;��-��h?����8���g�h��U+�\�
�؀�hssu���kF�_�X_�X�42�Վ½��nu��}�[�X�v�xݞ(�����S�����/���~@M}Ӫ{�������W�>���Y�2������U�qG�*�߀�w���'N���p[��4׳+1~��o�{��d$�;�Β����l��n�՝'����b��ƳC΄�����^�}T9�Z��~�z�h�v��<���(E~TYb�a�ĺ �eK
�!�K4�ה��Ƙ6R�n�����V����-tUQԏYZ�u�ϯAH�"+���0s�z����9���K/���������c����c��c~�V�\���ϰkص�)`kY5��nb����ǟ�VA��LG��l+���e�Y3��Y=�'�<��-b��nA��l�a{A� �*���7�*ւ��� �D�M��/E�uy�|l'+A��l"h�_�C_r�}���B�>>�T��UPn(�\ޗ�	�������]�3l�A��R�a��d���9HaA����A,��Zn���dA.�),��&bԫ�I��n����15�Zd�=�� �uH��,3�	� N�bD
���B������c��pʃd�`na����i!�&��A��%�����{�-�0�vAC�P�,�f�����&9ײ:��4X�A�ѕ,���L\����������X7�G�gY��؏Y�V��6�c�`��/)���_�%mXZ?֐���J{����#��gϚ��E���K��2��QB�zr-��%iX�U�.I�����@�;�<G��&]��z��4��P�l6+gt������&Ϯc��F�'X�6#U���zB��a	��b����(I�P�r��1S&RI���i�N@�L�<x��BOu�$�aG[ #!Eo����6��B��<���< n�s�y��?x����g�/�J4*O�~/@�e����������gr�^]B�Z�]�7�_�����P�X��A7�}��FY�K�����E ����k>�O�Kx�2��O���M�ݢĀ֫�3�K���|`s
�Cϡ|&{���;�=�x�3��%t�U�1W�C��oh�!��y���|,8׌��c�����؏����3]	k�B��a!�`Y? �XV��M�l%p�� Z�W�^+�|r%�3;��l�U���Y-K1��m2�I���p�W�aXͣ�������5���Ün�W�����c+Y=����,%��7��>R�Ah�	���f�6���mň�Y��ˊ 	h}�+�]�ǟ�h�~Dc���G�'�v�V�a�nvzO@ﾴ���4r�%��^{G�o�%@g"{�ƒrF�a��k'��cIߐ
�$O[io�ݏ���yI�N�I�J��;�M�|�ވ}'DW���H? ���B	Ԉ)�Z��"�I���r����m��2�-b�e���,�Y(��Y�Am�aƗ��G�^_��m<�m@����䰥�R����r�f@��X�{1�R�;p݁���H����sЧ�f��Y��� ��f���d��Y!�oA��z�Q�'����I�I����g����-��06	;�Aخ�8������3�DI0��u���F5|�B��ˏ�-�WX�VИ-r��}��?�e�ߌ�:�S����{-Z����r �D�W�<hY���G��R���[A�{\4����S��/��l$�G���@���C�{�Q��λ��|j/*�`��V��d��Ue��Q?w%�x���A5f<�j�aGC�Yv�����'�x@����d�M�惠�t�p�*� Ȅ�M���l�(FJA�x>�Q�5sQӝU�	����+��NE���Y�ȯ@�H.��z�t8OaE�>����@�t��L�BkI����:����0V$ET��Pr��o�5kEQ��!��o)�����\���D�TD��h�b�x��x�W/�H�"��"�,=3���U�){dl"#��$ǖ�Td�":+�� ��j�ֺټ�,��'��}�\�����/����uiU����������[3ZUs�9VK�g/a������[����\snDt]\���g����l�������\;6S�+�����Z�]�*���%ʅ��e���"�w��Ϳb��o��FJ>��7��}����a��cG����2����	t�A@^�XT���8��������"7x#V���7�0y���EQ�2~k��`;���l���6��X�o����!�Y������ r7`<��������*vJi�;
(@�xy����t\S��{�e<Dw\��o��`�g�3�y;��$�Yd�=��`I(��J[
?^�6�6���,b��t�sΈ���c�>�3��G����f8m���S�\�DVQ�·�,�~��R�'�d�bM������ھ���r�ѕi-��6��lǃ��pR$�B_tmOU���v�����
:qx U6>Gq�hW��a�y/X���A{&N�m�m����=�i�\�zXhg����n�ca}kώ=.������r�yd�gʂP���W��`��A��o��y?�P	�Z�IId�dB��S��j��v����g�S�(����r�}�H�.��bN�J��}Ly�3=x��;/���j�+{ȫ�Vβ<?HNn��1X)��f�'A�Q�ߕ_�#X�O�_�O��,������gX����R���X��"�J���yYo���}B��U�#x���u_���AI�����Y�j���.J��o���i�.����/ �*c��e��7�Ih�(U���cC�˼�v��R��t�M�8k�FZ ?;�<�����x��h��-�e�k�{�����nD���>�h���%����Ex�d�,Em/���p;v�î�=��� �T!����h3�MչX_�P� ��T��F��6��2ps�6K�
��ɸ%�Љ��j��Ė���p�.2AiNyl |�,���b�g��L�w�" �y&hAD7���81u�^5RF�`ȶ���Ȗ��(�A'�+0�C��Ґ&�d+z��ڼ	�l�>:��]��Cھ�_O��!h9��*�@s(�������vt6 �$�Ob���Y�pj��D
j��J�(��K|�#��dGA׏h}KR��T��:�%�2�-��'�KM��b-\^@�ċ���јWy���~H�jƌ�I#��e�қ5�t�
��@�����S�_��E��J�wɀr>��`wJ.�qw[�̓�K謐�����ʣ�� ��"��q��rI�|E��t�8 ��3|��)���K�#h�vm�.������`K��V�}�|�RW�r�Ȅ������]���
�C�Y�ay�Ñ?��B� q7�.1q����<�����y��S�~o)�¼�.;�/��_����38�<K|�W�C�AH�~�H�_���`�DǾ���h��Q�)/>f�|�����������!y�+�u�σ�1c�}2�&����{�U��߃��'��Į�Sv(��'�>������}��$'���� r�@��� 3<=��)]P.W�\�/c�uq(��r6b	/Vj-F�a=���W� ZX5U��U��B���g_m��=�����I��$y�m��HW�IFUH^�iHK�$#�Z;�f�$��S)��v�	i.�
;-�;����`:E\�����������i멱������&׾N�_��,��2ˆJ	��:��H��>�p�*�2\q�����9��������pd%;�v	K*�^ڂ�Z�"5ꠚ���7U��1���u���<�j��<��U +�P���<����R�`�AWU�뎸;�O�#�;a(;���n:j�'�O<)?'~qN~l�v�I��tq(K<�"�{���Ё��C�Ł�bW�)�������y'�����^S�}Z�������uꞟ�i{�=�����nS�4K��&��9]���	��Tw�$G�9]�$G��q��c��q��n�{ωm�ďL����a�hI�7�S|��M���mZ+�+A�;Qܵ1N�+Al�wV'kwf�;q��'��M���چ'ņu�m��j�-�e����[n���C��Y��"n4�z�[�%���U[�7t׷��q]����k�`M�X�$V�`�G�4�
S4:i�N�M��7�5����k�/I4�?�5���n�V���_��զju�E]��|�X��eO���`��A��X��R���H���'<��2E�)�k�S\���L�����0K,�E[�(*�|�E�o�yYb�)�˜Zy�(s��9�Zi��S��I%q��E�=ZQ������e��]��-����qNL?'���y]���"����$rb�YbJ��<)V�l�I�ڤX1�)&��Mh��9�����u�8�������+ƀ�1Ib��$m�,1jd�6*I�LY#��,���Ib����Dmx��$2Q��,�f�kC���G���h5cHg-#^dQ��ՆtC��q7X��Ǌ�G����j�,1��8K�H���T\Rg�P̀$�?A��N�R�D?�(���B�k���+A��S$�l�>h�'K�N�zv�z�"�F�ڳG�ֳ��i��#���#^��<�W�D�Y"�[D��"a��ʓ���D�,��şq����c+��kE,�b+D'��,gg�H��"�QC��,�,	��a��0ZյhM���}Hբ�v�����"��I����O���G�疻����6��Ӈ����~;�]ׂӼ�-b׊?�f R�(�H5x�٭��j��F"��D��$k+C�TC��'p���/����e�򒲉ak��MA4v �����BLu����9��s�D���)���c�xV)^��z-v�_q�ws�T��ɞc'�������~S��]�UlD}�#z��?$�sl���w�Dl�3�Q�Z٦<�.!�=N+��k�m섺��c��	�&�q��va/��j!;�^�mn $�'FkwY ���ڛ�d���%��$�pJc8���إ��a����`8\㤡��E��v#.t��نz��Gy�V��lر�F��㧎��5�_|j��~5*;����lqĞ�ү������'>�,N�{����Qq�_<�"h���b�p��Ay��Z�T�Ȅ�jc굠a��㢣�yk1z����zw�;������G�lg�CA+�ǩ�t2���g�G)Bq`%�p�G+
O�N��~�S��vA�#��9_�]�9�st/����LV���"�6e��㡘_:~��]<]cq�'���u��I��.z3���'������+j�����p��=�ųƔW<��{԰nܸ]������ǋ�"��<�䑇y���/;M~����uk@���r�+�>�k���Ώ��Ae؋���[���k_3�p���u��?TSյ8�gf��q'[�X#:�i�����]�{vM4�X}tOh-KN��3�Μ�;���ᩱ����Ǳ~Y���3y��[B�Ȭ1c�ԙ�*�V�]�����˲T�i۶Ms��?d�x7>~p�yf���{�?A����DXh��c�����Z��Y�P叽�7��*KT����}h
��F�a�NJn⻌�?�&F��%>��ȬDN����Dw>�|w��O��on2w�]}uC��W׉g������x�͇/6;�:rd��k�Z�Ք��Sav�[��;Y�M��k�j���$RS�n��ȌM앨��w����u*��q������W�W:��J�Wzi�������K�Ru���P����0?6Ǔ��O޵5�o�����J�ѻ�9v�`���x>���yf��7N���6�����
u������A={}����>]����,j��>ps���IO����.z�+=L�tw��Ik�C�Ւ���qz�������d�������ŋ��f�b?O�����C���_y݊!wW?��G���Jn�c�~���c��Ϳ}ޫ7�|��"��9�㸅���m*�.}=�f����nFL�&�YW6�T���q���t���IǤ1���/�
3��c��������+��<���T����O�Pv��g���gl�K�(�I4Em��rF��
���?^� �1��'b9�����)E�����^;��KN|�˛N�m�P	���~��;��U���j:��͟��%S$�Id͖�ĝ�Cj��r�8�X���ԮZU�lժ�ͼ�g�y��ӟ����������;���s�_��Ɍc�a�d���	�	":�%���ۍ�1����$;%��>~,�ZD���nr5u��弪7_?{�iI]�?��!���%�dd�LI�kh=�.9���Oo��~�;cd?˞��Pb�}���GLr����5ƙ�W���LX�T��oԚ��������}{9ؔ^��c�	)��a�?u�p|�끗���W��-�����lq�s�JzTztzL�3�H���uX°n�����'��Mw�7``��<��*ɼ[��?lژ�a���Qc��ޜ�**=o9�w��Ó�����^�t٬��������M�d�F�W�%�~������l�I��MJ钶kîC}��c���ue#���XD��X<�l�6�ĸ.�	Ҡa�Y������m��ms`q4Y����\_0��W�1?@���|�D��Y9'�{GQO�)�c�W�0��f��(�T��v9�\�&�f�3.vI6Bs���8�d��c��Eىv�
]�|�B��)1LB5�l���.У�{Es��^\]on7hn���.�z'^�XZz7�9�P��1c-m�v�htO���J�KS������"�{�1f���{M�יGͿ[v�$?��������k||R��7?�8���u�O	C����<�/���g�A�Ew</A(b�xA��&\��p.�e���2\��p.�e���2\��p.�e��'��2\�K=�I���e{5��[��pg����V^�n�r5"�1�5�y�ue��|�g߷�Nև�󝢿�޶�l����Ѹ;���s�r��y�E9g�y���Ո�ƒ�ev^gi��(�����w�	�G�|��iF/;�j��N�5���.�ir�Jwe>�U�ڕ[�h�{������LWN]��T�
�J���ד��]��쪪q7,�\n��U��jl����ry|��چP�2wC�5���s���<��@�����9r��@��ꡲ��S�k�pM`����q°a��h����U�j��7���4le���a���ƚ�a��Uކ�w��<I����^W��η2=��$Ȍ�i���.�rXo1C/�����5��0r-Xt5��o�ۿ���H%&��믯�vѺ���b��~wC�ד��Cxt���^����r7�v5b>��W��k�b�*0-[6�x�pWU���\6h��:KӮA)���t�܁���֍����zoC��I�S][�����Wݴ:OI'N��F���\�%2�ZV[���%�u��,U�5{$'+k�j|�M`���H��[��� �Kq2\�^���7P�1F�s���
x1h]Vm�;-��F��&[u4��_���4T7�0��:z|��/�h�\�j�%���`�R�*_��V��S�*w�o��$���A��	��J�4�Y�U�
Ը!T���؀�����k�]�]�>���b��V7z��(�b�}m�{��_���V�JCs�5���Q��C�[�����_�un?��j�6K�V7�d'i��*	�!~G�,�c)�]A��_��6�`��n�����C$�W����L@*S�Mh�xaw^K��>�'�J	��9v�"�n
��c{'���$�6c�+|�aƼ���j\��F,1we�WVX�r���q7�j�P�6���k�p��.��+��_I�$�������i��D�]u҃`��6�����B0�E�������n(8-�譫�L��wM+.*w�O+��S��*(s���+���s���>%�5��|F��rZ���/pOs�-p�*(��p�W��旕��K]�K
�QVP4�pn^A�tW.���
f��hy1u�I�Ib��K���mNnAaA��״��"Is��JrJ���-�)u��--).��<�-*(�V�Q�g�C�Z\���`���t*Ga���4'/vN��a1D.uQ�Lp	��y�sٌ��BWnAyYyi~�l�VjgzQ�l���Ey9��E��|���[�o�Q����p���Ι�_�6�lf�Ӧ�az~Q~iNa���$j��@���S˩%tM�S������Eڅ����ȧ! @�M%�H�"�+����Y�_P����)-(�,L+-�r>�C�8���Wd�+�H�]hh%{�����`�dザ���UU��&i����#�R�f��ZN &<��*�,�+�v�õ-.�%g��W�X7v#��zVx�ҕ`}��3YY���m��g�{wC�p+�Kw��l�_P���_�.+��Mp&.w3J��k��ooU%��t���4b��]�[���~��'����m�I}UMB>�ɵ��{ 8b�LW��|�W3?�eKY�gĪX:�Yl8`$r�h�b�h��H~楗e���5�}&r9�G�.V��;/�^�'����ay�-�y�-���*K��yI�*�����:�U��~��B�u�SFT$��hՀ$y���-$���,�1��mG!�?�{h�w�q��ޒ��ք��	�N�?S���W�}&��p��/�������&�^	��##�d�U�m�F���^��˦E��Sh�.�Y�?��s�?�\��r��k� �^�u��-������B{��?��WA��?aîo���֢���4�����(����)Y	ѫ'jm�kѮ�:�-�R����Ct���͚a��2�/q�@���a���&{�k�*,Y�lM�h6�W����Bm�!
���{];����a%)4snZ� ����m�g�`����4QMH?��G̖
��6����&����m:�%��>��L|�q�!	����KC��64�7��a��*p�LT,��$�!�dk���"%
����J��f�aF���|=�gh���o �3�A������K����,ڵ�V�����i��1l�M��M������4Bh5T��m�%�F��!,�Ƞk3�����m"��������=�q���Z��v/��=y��9��Em��4П�[�!Юmh�4^�D�s��n{�*�~;dk�6,O��|�hGr�s_OW�`�e���o5yI;���.�W�du��zZ}���CM��d{=����M/�j��H��_rK_͠�~!�<ĩ���m,�=�]8)�C�d=���訟�����<�,�Mst1.�I��:��b<f��^G�j/��������Ja��������w�v3����P����)a�;���C�nJ��Yk���>SI���k��B3���ј�ɚ�F�nX���<�7�#r�-�/�bj�ӻ��y��E}��X�]̇��f;���W�%㕔vs���ـ-�lIB�.��dQ�A�v��ɢ�/�g���h�c���᱾Y�J{�4��buXS��r�bV�;9N1���|ē�T'_t��C������P��O��8yI��^��i�K�P"i��^��B�"В}�Y��O/T�-K��l��o��=�k���^�3�Z��W9��O�bqZ��Q�sU@#�8���RПa��vѓ�g��d�(��4��ґ�,iNG�t'K��Z�ve����ⶈd��zK�|���	�����`l�B�<����#��-3HB)O���΢R��b{�e��J��K���:?lR~��N�_��r������t�0;lGsI��C1��KuR�R��ᖥ�2��%�Mr�G#�F�.*I�Z�ٹ�u�F�N�哦
�u������H֩�n-���[6Q�ݩ$���95߶��]{)�"�o��O��Y��ٳ;5<��deje>��|j�Cs]��4Z��m��FXXh���Y欽~C�(����Vh��3�G�ThsX�Ʒӵ|W>��*:�X����w���-*��?3X����,/<���wh�Vj�gk�j;�D�p۹B�d+�o�~Cч廭�Qd��8݊���?|��d%ն���i��ZD��4�%Y�ݣ#-+�tS� G\D��ڡ:�i��FYI�&;2��5�me���b�Sշ�AH�oӿ�滑Yg�ZҰ�'3m�~:���Dj��.��ì�Y��6�u�C��Fp�g��^M�c����������LaQL	�7��2f��Ma��Pnc\٠��m�6��U~���Z����ۘP7�� ���*򯩯#���>�'�0���y�)�?76�0�x��FR���19f;�>ez޴�r����+����:6e�߻��Թ}.����� ��$M�����S�A�0^V�K"���#\�W�(UP6��F�"\Hxvq!p����lT٬2�����|��zN#�Y��~�l�1��{����~�9ɒ3�%��l �v�wU����}��0��盭��u�}�.��w��Ɠ�[�IO�7KNaI˕e���>ꭄ�S]��!�ƒ�����Ԑ�	�oI�7���*��u�MdC�.�/I����9���e��A�#�AΞ�(�2��LaG����}l�\L
��
�烗j#�\��.�.�>t�ݺ.\�܋�Q���ӈQ��bP��,���׫롣$綮�GK�ˎ����/��~�����芡tQ��de�2X��Q&)���H)W*K�j�N�+��땛�;��J��]٥�U(��'���_+/*�+o+RN*�*_(_)�"�D�H=�K���%Ɖ)"O�%b�X$*E�hMb�X'n��U���>qPO�g���eq\�#��S�KqV���ƨqj��[MQ���(u���NS�R�B�J����FuV��X�w����ԝ�u���zD=�S_�*K}W�@�D=��Q�i�/�����%k���pm�6I��fhEZ��P[�Uku�_[�]�ݬݡm�Z���.m�v@;�=�=��Z{Q{]{[��vR�T�B�J;�+z��'�=u���g�Y�8}�����K�y�"�R���&}��N�Uߨoѷ�;���>��~XJV^Y?�������ҿ���Cu�8���ގ� G�c�c�#�1�Q�(uT8�rx�����0�O� ��5�d���5d��LX�2)X\\ƓZa�����:ء6��]��ֿ�	�%f��5{}�����V\��� <-?�|���^��w���j# �����C�A��jk�p������)ѡ��Y��Z�����ߵ���d�d�W�)���w��Ef#p}��k��V���h���$���ǔ���(�[3e����'���(�T+�SQ.$|e�^���픗%��SI9a��(³�d���x���	f���y����7��+	7��;��Cֶ����u;���p�fs��>9zD�c�4����D���:�JFɱL�bXYG|>�� 	+?f!�^0�Cyy���H[v�Y��h.��]�W>Ŝ����~��9���D�\l#�-�i�'a|_p9��\*�p�9KzA�&k�gԫ_�jI��[�Kb�w�1�J'�&�xi���|A�N������W����+/�_k����VD|5QXL�GTr_�?��9$�߃���o�m����Tb�?#1Jn�s�s+?9�|DDy*��������������#g������.f��E���^�Qj�C����}�k�,�s:07�I��7X,k�V���b*�.5F+�kJ������?�6�I'HW?��Z���W�c���H�`�Kk���גg�$K��$Z/O��?#�P�by�����^ʮ�4��x�(4b�Q��r]Iq���Y
bLi�7Ҙ�H72X��dLb+���=W6N��������d߷#��/�l�et�cn��M��%U�sJ�G��P�����-���>���՛ԛ�[���͛Ƭ�%�_�4)�Y�Е��3OJ����A�1�[���n�L��A���q�MEŀ�3�S����W%J�U���KIS2�,e�2E�Sf*%�<e�R��(J��FY�ܪlT�([��ne�rP9�<�<�<���W�Q�W>RN)_*gS�"FĉD�[��A"S�D��&
E��W	�X&�
q��Qlw�{�6�S���#�8*��ī�-��@|"N�3��T]5�.j���P���1�$5W�����Bu�Z�֩~u,�f�u�ڢnWw�{��!�	�i��������ԓ���W�yMѢ�X-A멹�4-C���iS�<m�V���i�Z�֠5ik�uڭ�Fm��Uۡ���i���Sڳ�����q��}�#���vV3uU����D�����3�Q�=[���z�~��ї��
�:�F}�~�~��Mߩ�����G���1��U�-�]����~F?�`�a8�8�Ɏ����1�I�\�G��ܱб�Q�s���;nv����hq���%��(�#���y^�giW���<Q���5��T���6x��<�_�}���S�n�������(Y� ~Tw �*0_�Jϖ�?'��)��ZW`�.G����]C�uY���L�eD4X��ץ��o	e�r�4U�<������b�Pr�T�)=d�Vܠ<ׁ����z O�����!�$V�T�9׋T�/�O����o!�M�<_Ix�\�K_��h�P��
�p�&�;��|�5�]�ɓT�&[&i+���p�Q&j/�����Gig��i/�rȨ&VG-wi���4D��)��~��]�C�<�'���u���*$?�E���LZ叨u��#j�,We$�k�<\~L�M�2B.V���&�L��5i5_�R��U����!��j���3��TrFbG��Z]��-�(�S*�X�ߦ��=Ң�^%c����dM�L�fH;Q�j�RK���j]�ܡ?J6&)�$�,�R2��7��d��mJRT��VGJ
�����&��<��=��Z�m���z'� �r��Lk��v�ܑǨ7��G�QZ�Zw_b��(��.K�'օ�*!O���r����I+��qD�!�*�G�����a0�1�3u�w���Z���^/�/�����ʘDW��x�*�
�S��ٟ�:Fa't���]rrR�퓫�}��B�r�?�!6Vb$��	m:�@7K��c�5	�J~�MFs��4S<��W�Wڒ.�i��J
5����>w�����H������]�nϐ�vH�BZ�����P��M4���+���7H�{Tɧ���.!-����a�pN"u��A�d��͔�)yԇB�TI��ٗ��?�K�xX�g@���l���4
g���|�ED
N;�Z��P5�"�k(�j�j�q���������8�S������2�W��Q�G�q=3��cxO�_J�3�(>�g�i����
~��e�������~7��o�;���?���������/�N�[c��7��Q�c�!���65�\X{!��\���Db��G#�K#�m�Ί,�.�;�_��w��ޑ�E����%lIji�������.�7�G�:��=/EYԾ@^�O<S��p-��x�c��`�o��]��A�=��}h���}��Zg�-��K�ɛ���-�_�� O#�~$�^�(�7�hn�Nl�|q3�sy.�@��=���_c��G�#6���ɦ`���e�s��UpFfSq�8��>,_���M��ݬX|_�ü�>��-ultld��M�Ml�c���1qkp�u�e>�>������A�wt>��C��X��M�[l���l�|#;=]a�\��F���EH�H5L�ʣ��.k��!݊�ic��;�v#��D:��ҳH�#������4��Y�zX;Y8��L�o��<��Zk ߭�m����A�Ð�Y��2;��aﳏ�)�<g�3���|{<�����7�����(�K��ғ���5�E˿��w)��|�X�j�����=�R����~�!.b��yH3�]�<¦�mӜɿNFL�,�RmD�Bԗ>xqlq`�q�c�8���}^��Yc=k�F�+�Yc%=k��xj���Q���9��^�g��E�N�_)rN�)w������9������@V��
zYIO +�	d%=���'��'�<̑U~:]�x�8O]�R6������jj��L�YI�����#����e�~ٲ���Sr���5=[�ԉv�ߡ��E�gZ�f��Bz�)gߺ�c]�B��Z����Yk,e��O)��:ߢg��	eS�ȧ������FĩS�l#��3�3�B��(5����J�ڨ1�uF��7Vk���[�;���-F����a�2������9�Ώ��:�r�6b݈5�IF��4z�� c��"��^�@��T?��-�7>3>��
�h�0��r��Xd,1<F��d�2�3�7���f�c����i�6�������3�O���g�_�e�	3z.#q�¢�E���z�z�w	�ȊZ�(�Y]>��N���T~�i�1ݘm��+���*�g��Ƶ��M�mƝ�&����{��?5�79�v�����/�8?7����ltu�^F_#��/��Y2�X�� �L1fRS0�v��� �5�X�`<��<�Q�l�a�)��Ts�j��6*=�r�P��X��C�B���&��_��8���w���'�zE^�x6=κ���&{�
endstream
endobj
30 0 obj
<<
/Filter /FlateDecode
/Length 281
>>
stream
H�\��j� �_e����n�B`IYȡ4�$:�
��1��}�	[���ϙ��3��}i���>�z���:�0�4�3�J���)���n[<έT���\���p�f�`�N�Sz��w��VkpF��uǐ起o��������W~;�_��f����F�b{���Bu
���V��?h$ɆQ�z�󬎆_�ɋd�G��('z"�D"
��g"JV�%�
]r��{Y�WR=N�J��)YY�F�ǖ�����saT�{Ҍ�t���Zc�*�_ Dg�
endstream
endobj
35 0 obj
<<
/Filter /FlateDecode
/Length 11013
/Length1 26648
/Type /Stream
>>
stream
x��}|Tչ���=I&�IHṓ��A��H^$�d&d �ę	!"�E�T�*6�(�G9�rz�Z��(Zѣ�Uk��X��G��r<-za��_k�LB@oϹ����2k���{�Zk2n�Q2.6�,�����gD�ΠutYI��Lx��i�K�j����'���򇲺%Ej�W=D�����꺼'���Q�6��:�o=���Y�icP���'�ۏ1O6w�k���� ���0��u�@E�)��u��ͺK?E���k[<.w̵t/����48��<<��<��-������W�:����z�w@o*xH�msm�HhQW`�M����<w+�wAf�����t5�׋���c��k+�;���RV�;�p���?�q�$>�?;�?C�3/�e�Q_��hɆ�`^T�>8^;����%�iE~lb���.��(��	����5�=R�ԙ��ѥl����MjV�1!�ù-V�}Lv����"ML�i.u�f�=����>XK��wߔ�_��.�Z�4����d��KR���X#xj��@����Jz�&�|�^� ��F/���%�F��q�2��Z�����Q�@��t�8͢a���ԟ��2�G]�ȢQ��+@i�c��NCoQ���z�VOoQ�)��o����^�<���`5z��g�G���f�q�|���^���J��R��=Fo�@e��L0��2��� �	G!���5H�h�t	�� �[L0�2t�^̳
��,��Kp�xN���"
�գ��+�eʻB6�c�/im�*6'�Pd��wi�������8� �{:��,�A��K�B/[�,�����lϰ�e��]B^X}�˅���t���TF��8������x���&`oR,"hm�xa9�����џ�G?���2ާJh�~�_�9�ǳ_���9�3?=DY@�_�J�;���|����!�H\��ԟ�@ya��,�JH��F�
Si21"���4�z�"�!
t�.��G��"���x��ܸ��[i�q��O�AÀ}h��̴��h-�b�0�FL����r�n�@��o)rD��4����^�]�)�"��R������]ZG=��N�x��&O�&�=z����n7�6~d<J��z*�~��D�i.2�j�^KI�7�v@�M��T���Mz�����I[�r��`ײ��*�{
<�a�٫���3�YY��d[�n�&;�X?I-�D��fo(*����W�ؗ�1����w�eˤ�l�0�������=���A�3��ؗ��&��]���ٽ(G@s������nb{Y.ke�����ͦ���2����+6�>�$��U�$3.]]�	�o�?��b�dGTE?��-e{a�}(/��CF/{��n,6�S�~z��Ը�f��+A����O�{f"ޅ/e�}
~w����c=��o��kP�K��.�m������p�^�)������M3�N���M4O���t����}��C^^H��m�)1�s�o���!g"��ۧ�7|�&�k��_͓��J�m&-��h8�K��]��7NB*�e�t2R&�4��O���������h�A��!A2���F�b-l5~��\
)���}l:�-7��)��r�#&ȅ�p���HzW��m�=�1��V�}��L�͌�R��|���R,����a:J?C��}T�!�m��ٚ�: ���� ��Ƌ#|C���(6D�p*��3�E_C7bl�̽�Ɵ�O_A�6�F�3�6^�M�ª�D�g�s���S�ht�#��j0�s�/(�k)Q��P&"k�n�b��:�`��J0� �<�݇}>X�Azc��#+a��kWs�o��#�~@v�S��W��U=_�B�� ���&r��h�:��i�Mo/Fm}�`ҙ�c	�����}vZ^�.G�Nx�j�7K�_�g�`٫i9�����W�
��iƭĞl&�W��pR��cn&�_�k!e�^`E^�0~G�#OM����? ��5}��ҧlKE�8E���c��ד�+dc�86�M@Fx��e�e���;��d6�9�M� �̒��x�1�+�B����7���n��l*fe�~%�^�w0 �=�鯘�`W�W7�e�ζ�?��R��F�C�X�\s�#B%b/��ˊ{>�)֦+����Z޿1�|�Q��*!��P����Y�
����p�܉���"��Z1��2��������dַ`���,"����55rwΏ��-H�&r�6`U�졽 �#�E����b��R:�>TD�Xm\'��0��ξ���H�"o �{Ƴg��}��Ǻj�2���\� j=r��z��k4�#��؉Xx�׍Hz��j�|B7 �������d�Ւ{1�:��`���ōr�7�x�@,˷�= �	���6�	L���eXIc��~)���Z�flG�M�հ��~����{
��C8���S���^p�݁��� �M`8b�*����/��36�/C<�7��㕝�3�ByE��`��8sUbm{��{�M4{bb.�IAVhD�e��^������s������	������!�(�-��9�
0�-��#N�1X��B��}��E'!^?�#�n�B�#�>!_�ܫ�n�_�QٸO�V���c����C�ς"�r@�O�Y=Yp�'��ŀhgT�*i�h��p�Dθ$\+��+���{"�DK:2i�ȦP$�﯃��Ѣd#"�	�Q�;��� ߱���N�ɯ{�)l>�'�
ᴈ��~n�|��0=�>����2�,~^X6�~�8��OKe1aYD�`h�t.l��Ճ�&�g��s��S�{<H�+��n0o5X	�t{��މX{HɦxQ����>�EʨZ-�Zо>cGno`$�������Z�#z<��u?ٍ����/[B�g��P(4�]JGh��d�	nLZ�x`g#$�+_�t�>B�%���8\�J,
��ٱ��0N(#؋8y\yWF�+{Q��c�~A���B|'�&�7�M!�C��e�u���q�h�l-�U.��̷�	���#��o�uK�-����k�9$V;��愨������8v���GP�D�Ͱ�)��
���
���QZf`���t�ǉm=%A���v�����wu��8���n� ��}��t��N���+��l:�N7�g���ӹ�!�+���q���;�]8�/�����S��b��
�F�f�a�,�/�L�V?{Mր9�?bď�bMƊ�)�K�鬏�.=�s�}(=�����W��c���H�9�m�]����˽���p�=����0b�L�s��FkqOA&��;vyR�}N3�#��p������a|0L
�|�����u��������W��˴��w�U�(�V���h�R�c񠔡�o)DD,BiG�@Y��G�DY�������X��o�.�1gr��s?N��}�}�B�2�-4	�+�틑o�H�k���_~��6��$GsT���7h/.Ϙ�3�QsFi��`|��g5�Q����<;��-;���u�?5gQM�v��k����5�*�Ќ�Ғ�ԧl+��m��Q�o%�?��M��q?��c���c[�����3�k��w:U�$�u�[������������Ο�������W[�3Oߢ>��g��=}d���-��m�#OMP�,�G
lOM�O�S�<���'t���/����?���@�1����
ۡ2��G���{��n�3�|d�zP珌���7����?IW��?I���'�u���Sտ���T��^�����:�y�z*�o�7��?����|��u���v�t�w:�si�z�h��4ޫ����;t������x�6�O�{���=:�U�u~��oF��:�n<��P��:�o��=˲�7߹㰺S�;n\��8�wl�ݸ=[�q����=�G�7��m��U���v�η��:7����&��cߤ�.�o�y�΃�58��?�_ӑ�^3�w$q���uަ���j��oX�T7���N�u��������q���sy�5��Fh�1���V]:_�f���0_�Ͷ��lu�*����Z�t��+��
�X�����PȗA]˲��$�D��:��MR�t^���F��:�J*R��x��+6�EWmQ���-�<�/��e:/�y�΋f�"�p/�?U-(��,0�����J'�B���2��ϫS�{�����yu|�$>G��|�i>�0���:���i:ϛ��%�\7��"��CN
��/���>I�mSՉ�|�γ���|�γt����dL��8>nl�:���&�1��|���.������G��t5_M��#�g�#t><:M���t���'��a:O���:Oڤ"��� ����T�y���t����ܡ�`��yt�����F�\�T5��0�6�s'WFsF�����Ys��ͦ��Д�G?���,���G/��g�e+a��[y	�3hy�^������><a���[������*��:kq�h����z�e��E�'�w��iw�lu'��IǎP�T��2�� ���Yi���.�������́��+S���cG�W�|�~\�;��h���De�ץ4�'�L�
�ճ|%�Ɩe���%�����U�8�ʢ=�f�m[+a�ľ��gOQ�lk�{
}ʿ�u3=/e$:�ԪUjdl��}�Ǻ��?ioSt�ж��G�f[�~ 3'�����G٬�6Z?@S�ݼ����+h�ݩ4+_���������x��-�>�Eﵵ���ǉ��q6����U��=w��tr;q�ĴaII�I-6:��|��F%|��}2)���Ф�1� AeKl�8���n���hN]~b�4��%�o}�����g�+SD!��ػ|��8R~��M!�m�c�͛'8��4���jG��/����a_Njh�ѡ�SX�¢�Dqզ�쪪�b�8�s`���R8Es��F!��;b��
���l����>�����K���,�����<�|�S���kY����G)��UR�X{i��(��vcN�9U�}X�3*-zdL�*Z5,c�`Y1,����X|;�!K��y�)z��AO@9qʩ�SԼ3�Q�_�����V��o�n-�Hr*����r����bP�D�)c3Ԭ�Y)Ô�d4d���g�g$SLO*�����sffV�=1#+y�=v��1Y ��I����'><u�y2i^��꟡Q��.�̞q�+��Y�2�Q	,5%�_�f�HKMQ�9a"�j�2������<��]3��oP��߼��څo_׸#s�/Y�/��X����m�V6,�Էy��_������.��-|z�>��C"�55��1񨤏PF�=MMMM���l%+YMIM��C=Y1=#=Y;�ݜ:,%-ў�2ܞ:&�;f�����	����`I����XH��!�6�e͑:�=+y�Ԋ�p����6{��6}nہ@��Zߨ¿w�豚�E/]纝��lي�۶�hX������������=,�u�eB��C�m�UheA&��X6ayVO��[�=i;�=�P�FOp�t-�9Q��<H6\�$�Щ�:�<9�`dKL��G>�S|��K������q�b�Xشl� �)������������r�N����d���_�=�#��[v�]{^�+{Ge97�<t���Ly��ۖ����LO�6+���牿�1��ɶ�I��"L������8������D�։�DX��%�)Iu:��9q��I��9�%8iDR|W�d'7��GY�>\X9ٌ�S'������yְK�\j�ëC�n�����aJ�e[��������i���X��W)��9�&.^��Cg{�)g��o���Z��8b���1O-sjl\l��"�E�������E���.��M(C�Ş�`8��i�	B�cωn�u���Ce0ȑ��S�d�`3����#�m̙�1��~�_؞��}��g����EJ��v�w~�$�s!���.)C���!����2lf�y��v�6�Ylk�������V@�XCIv�;�v�z���&��ce(�A�L%I�@rҬ	#��(J���;:P�<�r�U�����ojU�����_�p[ʢo�a��|W�����~��%\�$����Km-�crݞ����Y<%S���q��b�cxJJƝ�b��Qx��&���WiLJOҘ��Iv+�=�M�B�226�#�A��m2�;?��s�s`��50��9g!`پ>6�o�?u?�h��E��ֽ���;�N���Y濎�gmw�m���=�{���_�|�ʏ�ٺuECÇ��;���;
=$��R�c���î�D'����XTjLLt�.II�)ag��X�ᤨ�����d8�o���Q�='��������p�}S�*���	���T|��,0�w��|��ٷmk��t}v��� |g6x�L(�,!^I�S3��d�XU���c�[-c+l���V��$�z&�L�\��fč�b4:*1*j�%�ǞyF�G�Y	۩~�����о$A��`�����*X����.-e8�lb�Ĵy4��S9+I-I[N��re�d/y�W�N�n֭S�iݓŞ�.����q���F�HMd�K�K�M�Y����Ŋ%���2<m3��?g,Ԅ�8!ʛ=k<�f��UvO�����3��wr�����?����sɎ��Y�{����׼�q�MI�y�c�fe�=�ke�,O�ض���3�ף���CJ�����HAjz��X���q�X�mb��OQcS�.�v���62}Dj
�	Ն�^���4�����ۓ����ϝ����IFd$K.��2%#��9�D��t�����n�j~u̻?�':�K?>�M�R���잳����V4{�oczI��v�R���#[�m-d��`q�������qjbBʰd����SMD�L�vG�͏K�4�'��v'�'&�pg��4�%�$�q�GZ�k7+�}ƠT!�9�?
kZxQ6���/����˞��UK�����?�e�?��~g; 2ivɈ�%������}5��^?q��`�a(V��ol�O�U��ia����V8�.U��O��"\��p.�E��"\��p.�E��"\��~�?eLc	�߫���/P9�d�����/SG��mu��˪�)��[�hJ�����/[�z|�^��UO�Yh��l���G�XuFZl�UW(!v�U�4-�n���4"v�U�SNl�U����Y�Xʏ}ު��7ժ'PK��ž�n�w]KP��4Y�1m�L��[+�A��Ֆ���7�j���Z��j=��ǝ�(�w-�ԚZ\��<���h�v�����ۤ�}m.o{hL��=�U��}Z5z���,��^_�6#w�s�"FL�FX3�}� +-�`G~^��;s�N����_��m���y�v�gSnGKG^�����,��gB��Tڤ�ǣ5zZ}]�s�o!G���?��4sX{���8���A��`Q�]nO�˿A�5��p�x�mހT0F�x��Z�w�=����1C{9ZЧ�ڻ��|�A�m_*M`Z��x,C���|m.[���Դ6)S�$s2��5W �k�@l�l�]A�O��:�$0�	Z��9��gN���=~����#Ѹ�����HLȁ��Z;݂�.o���3m^���7U	�����hm)��o�%'�F�����k��^�j�?��`h;�����$��_۹��;�� ��>-������=MA�b�.)j򵻽B�@��Q�.W�o�GJ`z�d �� �0[�U:�=���-.�豴6��r���~����)����4�@(�dj`o��[�o��^�h�� \ u��RrSu"�\~�����KBnO���]������% &	u5I@��L��8��0Wk�AH�y!^�1����n�;��!��#�$ǊJ@(S�&"������w��p,f
ڡ-S�n�T�ce'��hX;a!�F�7̘gSQ��::b��V��0��A�iq�W =��r���:�"M�2�LS�Y6�k�-M'��ZEA��v��6��A0�"�}(|{�@
I,zZ�SK��U�Z]���e���Zy�VS[�����D�,��sf����~a��z#j��k��ª�ڢ��������N����+k*�K�V^U\�����L+¼��z�����H��TUyi�@VYZ[���E����s���U� -�j
k�ˋ�T�j5Kjk��J��h�ʫԂJie)� �����e�s0��9Z}maIiea��a5D���\p	Z�R1�naaE�VT^_W_[ZX)�
�UUW
-�*)�/��ҊJ!JaQE��D)�(,���J
+�J����a�8���J�Jk+r�����rQ��kK���H�����WWՕ.^����A�J���%gR�*�+��W�ևYYV^W��֖�	�V�]aO�2.�>��,~��D۹ށQb�%`Iia�	6��*����
߶��L�2���3Gz����e�\�MV�ψ,���?�Ē�c�_�>��X������A�T����d���H�2��ֽ���0+<
��Պi�0�*� v�������L4W'Z��k���o-U�%T���:�Ry7zZ�s1�/�3ɉ���6Kt���`~(��u��c���9��|�Zw�����Z(HM�&��������5b�FE� ��<�6�Ak9�c|.j��
Ш6�+ �<�{0g#�n�tP	j�A��E����1�#g�$~X�q���F��b���>�uɾ�x�$����Q4���^��|�쓸g��H<!,!S�H�Y�2%ZZ��W����t�m�߈����Y<r�_J�����KP�b�&�v g�*�<�?-���Y�v��J�YiO$��di��{�:��l�݅Z$�������AP�����7�쵴��~��j�������ċ��F�k���=���"�<�\�$�v�n��Y�z��L���#��I���+JL
>��#��^��,M��C8�����¨&�!�1��u�OkeFxI���KƂ�$_M���3}�	^�&�eOH?ͨ�Z~<)�c?�5�AĂ��b�NDK�>P�|�s���5��>y"�p~
9V,5��N���I���!��f�d[�D!��^ir�)u�aQo��ٺ?~��s9r�r��,�I�f<����VZ��R�4gr���� �뗨K��[QEC�̰햄��ny4r�]hb=F4I|�H?n��d�BM��[r�8͗�Yo��1�Of�~D�~��	�j��!0`l(V:����4)�˲Tc8o�|�Ԇ��]��O�H�e�6y��/X[���6�, p��ԅ�
�t��o��畱�h�������S�Sw��#�.�~	*��:��%�$rKN���#����*S
�P���wC4�'��2E�8� sI���9Ho�^��1ǲ{���@V�[�#�k�7�{f(n�"+�yX�KJ��3�X3�r�!ƇV��o3c�b�:�(���k�!K��sz�Иؓ��F�� ���KfVOxF��M�/1-2�k��x�H�:������Eo�����W��+�l���l@f�К�u��;����o���Cz�\�Y3�Esg?x��#c�_�F+F�ֺ���B*�t��K��j<��2�'ke�xA���\-z���%�.���|����e���򕈚��W�{9i�&���"��.1�T��EP��X�Q�+�Z�{�5N�/�Y�gQ/#�5�UaV��1O�brZ��~��*�C�U��Z���].�	�s��D�*����B�#�Y�,G�I�.����>��&�UR��7e)���09*�/�Z.G�׋�K.�zkd��P�S"���d��Y�eeQ�ǒk���C�i�r����I���-�m
�?�7�;eCe؏�H�
��%�"�'�(�YYa�b�/a7�y��T(5R7�$!l�3�w�(�I�J��*��:���b��"<_̬���8M�7}�"B��RFa�ŠZj�T���@)���KaZ�кG���U�u�ö��^v�V��X,��
����ZX ���|I��������0g���иo�;L\!�-X"����.��o�k�R�kM�c�k"�\�#w������g���ȝ�����ضA��[��l�Y�g��=�P+W�l���w��݇��ͳQ���-���^0ޕ��/�3钽�k�yl�#"�{Iה�Ӛ1���t�݂�B�Z��;�zoR����3�uZcE���N��A��o�AH�oҿ_ڻ��3�WjX�'s-�~
���u"4`~�6����'����}�����ݖ����M���2>G��V�_0�#���a�-,����C�<�6/1�z�z�6�ZQo�]��fG'1�FG)�M��c����k	��J��,����M��V���i���
�C1����έ��L�Q��-���Mޣ���R�(�FI�\K�h'�B�ӝ�C�O� =NOҳ�"�B����+���З�3s0'Kc�Y&�$�b��
�V�jY[��l=�`�u�;�&v+�����c��BM���vߠ�K��d=OOA�S�W��Y�&�7��Zپ@�ݲ~�9�����s�4���sx�L��۝�����s��3�Y�+#ڽ�=R��z$?e�>5��s�KTPW�Ti['}F��Eҳ%�\�R�rJ�R�[I��pL�	�w�fW1~�N�ֻہ�azl�ٺ���7̈́���H5Q�o�̶�v=����6���*�ү�O����s�_�a`��-�A([��^@�Ņ��x����ZVX�ky]�F��B^+���X%��/H�X���:�"qY�)[��yтxir<4���Ezo�5	��5G��z;^�wG"��L#�	7#N���țd=�أ���&�1�
���:RF�Bv���q����Q�#���C���v��<��o�x�Uq���N�>��?�Q7�
endstream
endobj
38 0 obj
<<
/Filter /FlateDecode
/Length 280
>>
stream
H�\��j�0�_e.����ۂ��/z�v &��b���gd$?�L�$3�����!�p�l�C��r8O���@�����D���(��u�86���,!��ٻOj���w��i3��Z������x���@az�M�َ�
y��c����Z-BJ��Ϙ�VHt�eF�%�
Ш�Pٺ^~G��MҘ$aI�$YNR�LL̞�8��L�$y�������������`�`~bʘ��SN��/�J�:�\����m��o?h'��h�
0 H��
endstream
endobj
39 0 obj
<<
/Filter /FlateDecode
/Length 1005
>>
stream
H��W;o�0��+4�;�� @�&C�ڂ�C��(�!��C�(�)�a��T8�δ,~���;>R83Jz�'��?0�����.�=���Z
��k^y���!��L0Bj�(֯�~�B��$��{����t?Џ��B�0N?�K)�J�o魥4���OӚQW���fO�<=�pу2�*�x4^�}�GF�"����{40�@=*V��{ #��l�� ��-H!�ȟ�չt�}����ݢX�߳7 [t'ZG�9;�!s� ���
��DD��}D4[o&F|d�,a��K}�`O�97Ƥ���U��G���#'��E�}����
�l˪��@��O�����Fal��~ɲ�w�PE("]Oh�Z&`��75< ��,Έ��J�nS�9ժ�mr�4�k�
�Ú���}���d��clu
����4��B]�$F���i|T�bKyB�;rF7���V��jj,y�B]�s"�YIO�iM�I�<��"S�2SQ閼�<�\.^������傫�����[�PI�C���ߢ� �����q�Q�SA�{��V�F��\��m�t��K��Z�5��/�ir�9V�丫u�X~���49n�srܷL&*�x�x̌V�dr�xwYȦ����E����M�0�P��9ٕ��|�)z+R���)�:p� Yg*�R���n��QCWS#]u���R/���e�:� �
W��'�hU�&�
�"���*6�m8Е�]�K����9����{W�*h��ݘ���7�m�M��h�E��z����Q��n�{�'霊JY�G���N;�oI�-�/@�C�*�����"�I���v`9�o�2x��ٮr�d}���6M=@!ߔz@��(KT�J����ww8P<$e��,>��L��|G��&�d�
ӱ2 �؅��Q��iV��iG`s#��X�B���=h�4y����$�p��;q0yA;i�V]r�����6�9l�����#��<��  ��.`
endstream
endobj
40 0 obj
<<
/Filter /FlateDecode
/Length 1054
>>
stream
H��WMo�0��W�<`�HQ_@Q ��nr�lð��i���8mM;�!H�Ȯ���H>~>������h����`M���� c�K��a�|c��o��F���XM����zr�߻z"�'}�'����u�ə�	���q�?NH�>�b�����oß�?�?|��0:
&�-L�L?�$���2 /����=�~ߙ�#M�"M��P��P����k9RO&���xHc��7����.�TpV��V:���-�N1ZCg)ʺ��^�s����hB���w�5��1A4t�.��v��0W�M��u�� �܅��:g�<�VH�2Rq�$�����9�u*�d�~�7'��.�>{�����m�HVZ{��[,�-%/��T��?�������TkVEXTj�&��fJ�<���kĔK]=��kP��	!�'�t�>#ڵ�h���~�D@���x�9O�(��:�Y�[F[1��-��i�+��6�'�X��]�FUl>�>��I��f$8+�����*�X��� ��p�V�`���8A+#�]�z���7]�X2�*{#;�m2k��#nA,"L޽C엩`|�؆�Ŵ/�eS�p��]�BܢЇ�h��Z
�I���$7��e�hr�i«��Q0�\����arP��U����Y��n�T��^7���{9J0�ɛ���v&c/s���c4}l4��E��aM��:Ĺ�_϶�\g7���)WE�+�� �܅��:'����4�)��k+[�@{ǃ{�<�������ͅ戋)m��k�K�e� QP��U'n����7��� �{��T�?T
XW�:�an���{XLA*ܖ�`\ҙ��qxՄ��*�9�`颎/�P,׭Z��m�����.�}E�Y��I�T�Щ)bwE�g��eA=>'6�4���(�ׁܢ���`J�� ]��N���A��v�����w�ir�-�̣��hI[Y�x���y8��u_�d�^��R��S�s���9$gj��L>C��`
S�y���Y�,�|!�u�@�Ar�ՙ�Y�D��Ř��  F�3�
endstream
endobj
41 0 obj
<<
/Filter /FlateDecode
/Length 1005
>>
stream
H��W�nS1�߯�k�{��P�&��Rvb�T����f�֏�U���;q�������)���	�+�q��_�O��i���U��f�|����Vz���<�>Wkt+D%l�����SY!��9��<�[��kt�Ѕ�P�N.�V�^�J���:#�[��}Ǆg1��ӌ-�h��0s�:�4N[㍖��!���8���ÿ=~����|�z����[��(aL�}/B����y�o^9G���1J}{�̀�"hzKstA!)��f��r��1jA�h/!���pShtR�>ӗ��Ӆ���Mh��P�y\z'4\�:Az�:7��`���#8��i�.�8(-T�� �*`��aw�5��$X��V2��bL)�mz�Ōh��k6M?mR��8����NXwu�m��������j���F�s"f��WlH�gh�I�֏4 5Z`��f���;�]9@}�����������>ت1cMK�qdHφ�Y	���{��5"��=t�]����eYǒW�S��]�� �Og����H3i�(o�,^/IjE�1��f�MP�ɳ�Fr�g�=��wl��"�W��Yf�8T�S~�	^�������r�Q�x-��K�ѴV�M+B�l4E��r�0�&ko5�4z#z�|�̮4��͖���S"SYȢ�^t2���l3�:F�g$G�~�h�UAZ]֟M5X�����/0`A�Q~�f[!�)ԃ�dh�h��Y���!�ĬB�wT2凞�����32�_l�=\��e]�IO��~��90\���9�ff�� ��4(b��f�U�l,�Ԑ�<X���S��R����n��n���ҢG8�e�h�����.e��):�\cĉ��w�����i6�y�����xM��O���tc������Q9|]]�٫��c�ʬ�(��Y�*��_�`wɛ��Zm	�U��yp�hro�*{u�G�I$��y�b"�N*�I2H���	�Т���j�jsj������� ��7r
endstream
endobj
42 0 obj
<<
/Filter /FlateDecode
/Length 775
>>
stream
H��W=��0��+<8���/��K�t+���T�-�p��CI9�H���%�T�H�(�����H��e�*�� ��/�����x<����Mq
x�G��э��� ���4�����܇k��]���=���#�WD�qN�t$���@���q#!��Q�?<�#��_�䗗_ϟ�ߌ#Eaq3覠��·���&��b��%\KJS	��P�p�	�Uq���z&8fj�S�
�j&�����]�\��.�mM����f���?]�@�3a��@�E�U0+iO��e�T���\sl&��
�Ը����Q�y\C@���Q��Zۜ)����,=
^$,o�©I�%Z����5E��g{U�r�������k�t�h����ZȒ\^�ĥZ,�:�F�Yhv�	�V�Ǒ����McI�+�X��c.V�.������fq���$y,�%�C���q���֝c��W��$��j�-�c��U�>����/�-�H��M���͗��.�� �[Yy��dSG�ܩn�����:�ǫ߷�<�!��	�w�E����_�_��s`z�/�.�u�N�ΈF�o���eObm��U�אq��n8�m��j�y�z�h�Y�m�Qb��t�c�)�rV��c����dչ�<ЁU7���li��K�Hd���*�'1��$'OMiFvɤL	ZMW��vj��V�)i����-�`Pѕ�㩆u2F.1����y��;F��Ke���'��	��{�=��G� �)�
endstream
endobj
43 0 obj
<<
/Filter /FlateDecode
/Length 665
>>
stream
H��WMk�0��W�\��F�CYhh.�|+=�R����:�D����Ƨ�k����=끶*bo���?v�y������J�S�Up���n�����|���=э�7=Z��hG�gx�����).��'�	x6�G�*�03����>N@�hjB�_��A �<0���Qk�.wQѽ���}��=���h (�M'�i�#)FN���ii���������n��
7�Y�sn����m
DQ��V��y�S���>1�p�j+�v*l���W0]��Y�CeEXc�N�Q-��Es��/��f�*�NgJg���؛�b��TU�{T�,`���|� ��X�<�K��pKЮ��<Q�G	-�=m�M?�����R݈4���l����$����R'z�`��t�����#�������hyi$F*Gܶ�@*9u&ZE�0U���j=Ep
�Kj�Tk�|κy�a����k�;���!8Å�u��!i}�<��#ܫṭ[B���C�vޡ�X��Chgyqe�G8�����;O�8�LA�&�C�{Ѭ!+��Ch�r�!���:�&��u�n��X]� ��Cl��!�� A� F��H\Bٚ�8�7Te�tuⒺ:���z��<;�!0�5S��b�C(�<��y�m�� x�*
endstream
endobj
44 0 obj
<<
/Filter /FlateDecode
/Length 736
>>
stream
H��WMk�0��W�\�зd(	�%��o��B[J����Cglٖdm�+�{IX������͇�{׎3gz���r�쿟;������~�:���)�kc�`�<}�c\��%�������~u?>A���a��M!5�xZs&}?��Ϝsuw����fz�M	D���U�
mz<5è8�į��ܟ�<�\��G?��F���O7oAr�ܞ_��Lﴸ�^؁�L��,�b����x!3��������D�BB�؝�C_��S��Q�H1��dA�pX?�WWҒ ���y�Kq)�*\Ah�Fe
TYf5�J��l�m~�ش�����'bV��c��Q�j-�A��������Y_���u$���.�'�+������9���*�CW�a�ԕ��X]=O�4�~�*���k�� l*�35k*�X�������RI�<FC��d��ڪIIUճ���њ�#ֻ�uѠ���NbT��dk�C}I��Δ42I��;�q�^D
��M�dDZ�\�[c� �������h$nq���h;��p��a2�V&�۠*�`5"�B�3h�&����0�<�^\������-hG�b,V�뵻�D���=Ө���v/���&��<Z~�{��.����[�}��P�'�w����@'��Y*?Gx��O�����%@����2�}���O��YD�J��@eQ��������Q4 ��8���l ��	�f0+���  ��3K
endstream
endobj
45 0 obj
<<
/Filter /FlateDecode
/Length 719
>>
stream
H��M��0���>vЌ>%д{魐[�Ж�9l���#��Z��!��`�������h���Q)��{
����!��~��=��N�����in�����x��ս�->�^� dz<(߉ݧ�C0�x�h��~vn��~v���ނ�
\�z��NKSzw�s���@�B��Fec�2��_�� ���[�=F�v�+�鬃��b�!T���/��`p�����u��U���s4���UqFu�a���81�Ժ!�x�F90�<����~�d!yХL3�]�9��y���pEJ#�i����7`
m�ⱎ���U˪�ZA�V���XyfϿ�谸i)���K��&ZZ�eB��J�f��Q�Y�S�W�t��q{�;t���ul�ш��O� 2'�n4ī2�)�'��1l[�km�L�j�H��I�ն��G��PkV7��n�X�j�6Wyy{IW��oH��(�;%S�c�ae	A�ęL��H�&��kV�n!ȗ�3!,]�N�H�	!SGz��n�>WB&��)��ýGoi]K�69BHW^SB�� F.τ�+l@���^U�@kB��Hs2��F3B:��Pa�!�x&����FY�hIb�N� ��L��9Bv$1'B�0q&�<5[µ�k��JB/�3!$�o'M�+�	!SI�w\��+�%`!d2[�2��1ܻ�pI�ZBȴ	B��B69B���'� ��-�
endstream
endobj
46 0 obj
<<
/Filter /FlateDecode
/Length 884
>>
stream
H��W�n�0���� ��Fӡ[oE�mQ�C��C�(9!)%N���ϒ�{|�{�t�Z����p��5��(L0��f�׿��#}�y3��
GoA�K��epAiG��ϟt��~��u:��OiS`P+m�*��|���p��Jk3򏠵;e\����x�q����PBt��祤��J��J&�\̖r����TC$(�9zd��Q+�Ag����cla�J�f��t��e�k��l��4�E��魈O����Ӂ�]��Dٚі�tT���s^�ZF�C�c?
I0v��;6�r"bSQrp�7Dw���!@俕�j��jO���"�'�6�]M��ԕ��{	���<�C����&�O	\c��֠"��q�m��n'�)!)K	�M�(��#�+�V�m���y��
c|L
SB#O��̑hN3S���,]��Ё +��Z�B�a"�ȍׁ�I+E;~�V�g�hͻݹ4�擆lP�zڟc���c�Lc���u�J�(�H��J-�ԫ�T0����t=�-\��W�}*2VZi5�_�Vd������X�b�j_ڟ���m�9ϷKj9!֒�}	[LuA�.� � ӓ�`�T�*7���&S�i4���M��&���l�ay�uUh�h2f��,ߢ��ej����u�E�pw�������v6�
�w*λ>G"fgG(�%�ʈ��)3u�E�����*\��k�lPV[$�e�*�^�ыdUm��A����d����J�h ��R�6��D�I��f�N��9��&��Jk�=�c���r7��n �aw�0c����>槩6f7��JF}5���ј�F+�C��H�l!�r��j���U*��ԩ�S�]���g:��e�� �+
endstream
endobj
5 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 6 0 R
/C2_0 15 0 R
/C2_1 23 0 R
/C2_2 31 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents [39 0 R 40 0 R 41 0 R 42 0 R 43 0 R 44 0 R 45 0 R 46 0 R]
/Parent 2 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [5 0 R]
/Count 1
>>
endobj
50 0 obj
<<
/Count 1
/First 47 0 R
/Last 47 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/StructTreeRoot 3 0 R
/Outlines 50 0 R
>>
endobj
49 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227153517Z)
>>
endobj
10 0 obj
<<
/Type /ObjStm
/N 25
/First 190
/Filter /FlateDecode
/Length 3735
>>
stream
x�ŚkoG���W��D���[�� @@�l��]V��g�%��9����S5'6�lm�񙚾w�[�nϰ�C�a��{��ZCӫ��n������ޱ������gPQO��TB�Uo}�6Bjz���[��X��r�3��Sy���9�FYb�Mo��]C�a�RCa.��]����������˳��'/v�����Ϗ��߽<{��|>����ǝJ����ͫ�k���ݻ�����|�1���z���nbC����ǻ��?�ňxt�`�M��?zu��mh".����_�'�w�\�V<�!O�����WZ�7g�g��ˋϷ��W;q8�|�����.?����_���������Ko�t��?�)������+/|�+-���d������v�������?��û7��l�����Bc�k�e������ow4��R�ֻ�����/��=<x��ޟ|Y�ӟ��"ԛ&�轅?��
D�`$��8NB	�^�k�FL)�h�4�)ֲ�٠���V����
��g�aB�Zk��s4kmJ�`�a!�
�����R߂}�y����΂$Ӆ�&�^B��]P�K�KU���t�:��j\�r����T�&��2iNa��*m��MZ�j��bDU��4��,M�R��u��֤P��%�4���mL�M�Zc�{b�'T�
������͐i]
�d��ԑ��u�-,Z�����X��51 ,C-�����ᴑ(�&�X��	�Q]��.Z=��n�+HD��5�I�t��c��&q�?���+s	o}�o,V֗�����$�kk�!�,Q�,�> [�8� �
oc#l�ɋ$ ���a ��_(9���1x�WZ4��"��n�@��t�"���`���UxP�ؘ��i�c��XAE2A".(^��`c����g�-�/u�*�;�E� w� lЀ��E{MeU�h���Q�L�(imh������B ŦC�y,�5SC������%���kHYoL`�)H��Z;�����k�j���R$�2PJq��MF���UV��֬#�\��\�G��K5V�kU]ɥ:����S�W��ߚއ�m�j�1�����fX@ ���ҫntd-k�qA�0���	L�@k�ʤRe3���\b��yd����.�3Ι�*_d��Է�P:�|X;Ù6R{q v��I�wY")�[H�W,A��Z����U�V�Z�.�b�V��f͂�Z�@��h@v���WSe���Kq�/�[氈�E�%���E��-��k}1�
��f�bz���p��Zص��\��z�ۑF���l�����bic���x_���A=�z$�0��N��b�>�.��h#RݚZUt��WNLje�Ke�D����u2_�.
��5%����i�V��CG�E�`/�k[�#�c��.�ͦd�"r0�����*�NA���(�	ʕ�JD��9�,F&flX�b����u����bCe�-tA��fpl"��('b�4�9�Wk3�xv�Y��m�X*8�Y�U"\��0uq����[pr�/��aɴ�rM񾉇�ib��Q�9%b��I�'�OntpU`O5	sR<�I��f��3o�[X;�k�MR�R��ۢ ����"!I�m+o��*'���M�3���J7}l��W!�&��C��$ڵ��`����VͧJն�%�(8�m)�0�#Pa��R
�;«����c^Y��{���f��`��͌M���b1F��l���I���}����dfX�F�����.Ad������#���nt�h�fG<r[�,�i'���]��C�ۄ�J5��Q��W
km�9w����8L����XE�2�Jt�d���l�yRi��Ǖv���]@_0��9���/���6��OZ�CF���"��CUM/��5d��<lG�\��A��|6�(��b���
�겑�h�Z����pcXnA0R�=-n`4�m?#�4��C�A��	��.��ތ3��X\l^�,Ї��sq{��`}�i��CF���Fxf����{	���L�f�a0H�b��:�,tJe��u�̭�j��Ӧ!9qc�gC1�<i��RC|�K�������ۃ>+��#�d�)�21"���;Q���MAn_�����s��}��lS��d?Z�4Xm�ې6N4�b�u?0zqf��ʴu3l% �$GĠ2>S�]�7nh�����Xn6&vw����-��_�����"u��#(�l��~���[��7k�m=�݂�n�!�d�wq#W�����-�K��$��vM�P�YQ� S�U$p�*��9��b?ÆA0��]�`�V�9?��-������fa���f�_.�$an�f0����~�6��23�����d����f {�1n��^$�����l-3����$��B����T�/�!�M�s�EXq3�ɠ����X�Ev�"'Kd��G`�$����r���1�0�������5���S��IѼ.:������p�s+�q������^"���k��	���_�%�f1J���0T�Y�~�0�$ �X��'�m!���ńRN��#�*��Y�ιH޲Y�'�׆yƅ�=֙�g;8"�%4���+�C`�����KS�f� �4b��eV�`��P�4�{hB��6-��ҍɑB�����#��7O4����ꮟM����5�&��r�H=܈ZN&��o9R�#��K�;D�@��Qd�=[�F�Ln��\9�ق/�^���aSF�Z$@�֒4-�i���3��1�'��$\�Ա#��~��Q���S8��d?\��V#4�B����iZ��ґ����l���X�jò���I�m� � ;<��D�3�
'!F3`v\�u#�[�[���#�&~<
�do�S7�([PI�"��qޒ5�#�G?�������q^��	鐌}�E;�!��w�r�_¿�b��E0������0b���G��[���e]F�j$�*��ܜ�X$�2�T��Wi��ND䧘#�9��������ѓ��v�yU$m2�7E�͘�`n������|xr�A]f�ĎK�v��6�Й'��<1�X�=����<R�NmZ�Nl�v���h�vr�M�:8�?��7
~����|O˷�������/��9>���y|�&�p�p��35�I�ߵK-�����Bh��=�ñ���D��V���~F��1�.nܠ�%T�k2���I��T��2({��l�)��*�Q��9�M�S��(.=�'�r*�e�Q�95B��
8�7�3@�_���oޮp:�r
�wj�@�zh�5���(m�#�c���<F�cY�S)N�;E^�g�F	v���ZN�c.�)n��<F5��`�<FM���cʆQ7ѽ�k}�(~������_��w�)l��ό�p���u&��p���ߜ��ҕ���z���5�׮9����궒�K������;��e�4↊^��d+�'L7�	�_*޽{�����������
��X?�o\��K�\*7 'k�.���K�V��� 7��������W��7����>b/�6~��
����?	��n�-�n�܄[���-�������������4}�Å8���F�>�?�������{���6�����W���탇߇Ϗ��;���u��x�_9��
endstream
endobj
51 0 obj
<<
/Size 52
/Root 1 0 R
/Info 49 0 R
/ID [<A96308C1E407714EAD36CD4292AB91CA> <3D12B16FD98D0B7B5B843F21ECB4A778>]
/Type /XRef
/W [1 2 2]
/Filter /FlateDecode
/Index [0 52]
/Length 166
>>
stream
x�%�;
�`������zO�Xz	��J��{�Y���� )M����v�f���q��X�Lt<��s/�H$q�CEn �F�+��v�I@*2+BR�tk�Ej�N��V4I�ubq@ڤC��|��>��<�)��rf�,��C�����#{6"C+�*?=�-�#`
endstream
endobj
startxref
64226
%%EOF
