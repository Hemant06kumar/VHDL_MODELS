%PDF-1.7
%����
10 0 obj
<<
/Filter /FlateDecode
/Length 22
>>
stream
H�:��*����`�t@� �+
endstream
endobj
11 0 obj
<<
/Filter /FlateDecode
/Length 3482
/Subtype /CIDFontType0C
>>
stream
H�|�{PS��o��il7��&�ũ�`y��*t)OE`uU|�$Jx�j^"�"�+$��<���"(B][q�j]ݕբ�V�]�X�����ދ�3��L����;�������Ι�B�f!,ka\d�'���J��P%������YR5�\E
�E�\��Ez{�"��:Oy���<�.%��#~FFq�-�m�� :#�"<���x��د��+TZ�6/�8��VL�J������538�!3�'Y���?�kf4P2�K����*25�h��P"�R�B�J�)#C2�Z#Q+4
u63�~;�F�PjSj��vT��j�\�UK�L�:]B0��2��R�JB�|�R2V���H�*�j:1SEFd��j�B�judRr�!�$T"W�_�4(�|� �9�d)�,���@�U� �� �(� ����$��L��z+���!Y�XY���bg���ك^Q^�9~�Qtz, �����ξ;�='k���%s�sos�K/��/�h���&-�<�% 2tZ$�6Pvj�sH�sY��A��0��(�"��I[<��W�Av�^�aA�8������L��8� ��rc�0->ƹp�Ҽ�@���ot�"}����l2F
�|I_�-���QK1:#@t�)��`���z��	��m��÷�^`�(O��^e�yu�l�~'8��ܼ�y�7}�]UF��̸�HV�-�S~�"pj�s_8r'�¹���%9���,Q�\�r ,4Z�Q�go �����(v�vן��:�6���C/6D�Ղt�6MyR�v��vwiN���<��֓=nM[z�F��ڪu�y0���IA�	.��a4{:h��T:�'caxL��3�ޔ�Ӓ��S�~!3]`�M_�r�9P?pb�J�esӧN�S�7�0�.��w?sO2`]i/9�͂�Ir�� �T3�K�p�2l0�h�� ��K��Wⱑ�/ �J}�sXt=~e;�R�|}5�6����: �3�S���]�S�A������Pě*uݰ������	����M:a��P��<���"w������!n�<��"��N��B�
͆ �J���*/?-z���0f׉�Y�Yi�����n�ID�=��h����`��9@�l����MSU]�
M��[~\�A�5YL�
�C�[��'���`H��A�:���m.�_e���a�;�R�k���	4��D�/�A���tV�w�k{�b N�벫r�2������b�MM��3�+TG��B͡8LM�`��n}h��Z��%!�g91�g��p�0����)*�����x���2X���r&~�&�A�.�%�7�����EY��X��Ǧ�J��@��j�{1���坭��sQ ��P���C��K��DO-(����o���S�Ҝ��F���@�Mc;6|�\��q�?V�r�Q����4��Br*�
�_ْ�Z�B���G{�t�F���O��J�L`�i�+��jҚ�BJ�!̗��qK)�Jv%u�'e�Ϟ�7�E*c�.g�={��\ol�c�6��_�x�=����x}����ﻯ�=k��m�`��+�#�4w��I?{zCZO���ͺ*9V�Q!]���=��~�
�`.�����=�G4� �� �l����"兑���;���#7&��	xU~��Cd�?Y7ZI�8�=s\O���PG��}�k���#m����v=H~�<y�]�Ps'�m�zc���<�1X��{���%��{G1�v�h{�c�F{��C]�@LO�Ц�!�Ԣ����B��(L4�-�s�(������z�����bpc���4�>�n��F��V��c���	��9���Nx$�~P7���������LG�0�(FN�`��EGqm{NC]��D��~���tb����&����<��~hK��{8c'�ۄ/N��8'��*p`�5��za�w�ܼ�#��c��˽-�}�������׭;K���9��`�s6�#��p�ps~��~	n��M��w��ϋ��p���/���W���1_�6FP�ර�O�ES(�m�U�x[Yf��	+q���y����7ì���!�l���i�}�$��P��ȕ�==��)��a�X�5--�5Ga�ؙ��	�[�e��Q�a�jc���p;R�Lu�v?n�������1�0G&X~+�=>�E���BY?hKm�Pz)���ł�b�!~�ЂH��(*E3tb0Q����嘸����y��}�s�#,��G�E�����Q>{B1S���+��E�d+�@�{F�9�41e�5�7kZ�����=r��B��Z�s�-�T��xpdC&$`�۸��~s������l��~���|p�WV%���&A���?vv��H/�Π+K뇙�A��$�Z��+��v�\��h�9L���������}-L+�����T��!���`��38Ç1`�{�L��h�je��R)�G�����,��G��A�o̕`�%���6�X�K��.I˯ �>$ڢ1��`0���WK�0�\�a�z��uZ���ЩZ�� U��lm��-&K��С��w���'
u"ّci��	��4��%[�Ɓp������/��@��(�x���x�+�`ER�T"{)Ҧk3���r�����b��04�׬���W/=ZQ 7�Lu�����ڧD��d�G�RT.W�J��'�A}ŀ��+�v��	l%�Xd�rd].��i#��v���[\�
>�`���Y�R��tyH�*7<���S��sDJ���y��Q��>�K���U}�W���[�;02�u��t�We;��K���F#}�7gq� �x��������ʫ$%�U�$�~��A����BreY?�7�y��25%�0I�h�{��a���o���4ԟ�bͷp�-"V$�	�4fFg�'��K���=Zc�$�	�� ��r��f]3M���<t-��B!+�c*�$r�]@r�Y�L5=�*�>	��@�K��))� ��Z�=
�3��;ǻݛO�o�xM��5F�b�"������H*��%ܸ�!��G`�k�� ���U1��ŭ0nN�Nޙ�p k��M������|�`M86���u &�Y���hD%H���I�&N�M^�p��5�hC0/HB��Oxx�v��F`�f-ihoA����}g�*�#i�[��Y�{�y��O9�؃Zj��|��}�w��^|���R����ޗ3yKƯбDdBk_���-,^|>���5H�t�\���g/�)���g�E ��3�覍��jK�P���Uw>"@�?H{�ɭnC!lm8�(`�e#k�9GC��̐�f��g3��x��r�� =�����ܲ������Wp���?*�MB=ݼ�*s�A6 ��"9����g��t�x�4�Ǭ��Lm��ɀ��)��d�o�w[^>�������@�G�Z��J�m�e�~�)b�g�M�,���ح6�a��YCa��w�7�3��8���7R��� ��
endstream
endobj
12 0 obj
<<
/Filter /FlateDecode
/Length 313
>>
stream
H�\�͊�0�O1��P�֏D(�<���l2vk1=��gJ6�G�τ��؜�=�7�=��(��xw�7m�$����r�l$B��'�Cc�1�*�aq�n��A�W\G��)t��`u9�k����x���Aaz��[7 �mֵ�7!��k�)9���Q�d;��37��8��su�F�[Ov���s�=	��8��EiI�
֞�#m3R�e�����"amY)�s�2�Pp�p4�dX{։ud�Y/�<f�Y\��z9�+�^� )c�˜����Ҧ��|yw.������t\|�v�Rˌ~ 9��
endstream
endobj
17 0 obj
<<
/Filter /FlateDecode
/Length 22917
/Length1 50064
/Type /Stream
>>
stream
x��	|TE�7\u���K:I'$��$MBXC�Y��!�$@XB�6Y��-

@F���A���,
�

ꠣ��#NTFLn��{;�\�����~���unݺU��V�Nu�nB	!�@2q$%e��x��BNV�����Ĥ��V���G���6&#�q�,!��"d��c�'�Z�(!G���%<���_����d\Nqvٵ�o4�*"�=�3��q��d#��%B����œ�?&ā6�gF6�2��:��f�͏�J>DHw���Nyٹ&'A���
�`��П��SAq�d{�ڸm;��4'����[�$w�}nq��2����:8J�����J"!9ո\VZQ�\B&a���yYy^Y�k�A�QK���Е4�6�_o�M��=	6�z�D�]ןV5P�y n����q�b�tt�UN?娠���y�g/E�����l���WА/ҵDAKoen��+{��K��Z�Y�$����m���|`Z~b.�%�S����fS1�l�;?_$�UI���(�HJv��N&;I]Gs�u�O��[d#Y���W��d�Nב,7I;�����4��W����=2�Uh����$��#\G�迅�E��D2R��W�I2pR����#�@�$�%+�Lr�$��)��u�7h�o����j�	C�kt((z���}�`��x�D?���{5�<��9�^����i�`2�`����G�{t3��߀�BdA'(�d�����F�{Y	:f��w)�-
���$�eq:����!����f�k*�[Ш����$d]�XF/�6XC�Zh��D�6���ޭ�W��w��*'������A�5�L��f��=Y!<g%�^}H{'�Q"<��� �T����6�n�Y��XH2�l&>�j�-`!�o�3�� %F�����3ލ�y�V"����Fqj�D�`�C�ǌ�]cV;lX�5n%-u����B�WXtV���ǻ[���md&F��s��"�?V�e��;�9�8t0���k�"��}=�	����;'��rZ�!� f��d-fM$��7��Lp����f��K�����⍒]?�'���0�\ļ�@�V��$T�v���(����,'��`�5��4�|N7�QЙ��onЏS �h7���8�φ�4R�t�A�i����$�1�. ���h�����|�P�6�f�nGަ��������a=O+��m:���~���i�����MΙ+(�E�$f�+z�F|"�Yr�A�ϹIA�V���Řo(	�ם��W�`�_�2直�������p8+<b���U"�>X/��:8�z,~c{�V�����x�A[I@��lGk��@[�3�L�=�Ĩ�b��
��H��@�N>�j�4�?!��#�	h���v�Yܭo��X\W��y��:_��ίHZ8�!�N!_G���\.4\��=���C�4ܗ#z8�q�EI��YH.R
��O��R���\'w�`|�.@}!���K%��*	���XK�Şd�P�8)z9Л�����\�ꍙ�Fyl&���@�ǃH�F&�����v��]'�A}�Y����<Q\t��V��ЫOM�)r~�D�9ч�f����4��b�w�@�:dASq��2-�@a�x�z\���~o����.�G>�s��#�/�d�`�[���z��!/�?��VR�P���2�#v�S^Fl(@�ߓ�:���ԉݻ`"VŻ�C�%W�~J��$%P�!}��hd!_�/��� v�����s��dyR|�b%�AV8�&c5n�.�E���`;9C�a�'1k��f�9����?O�P�1��!Ed.r�$�T��O��3�()s y ;���y)|�V��p�O����_%: ��!���,4�&;o`�m��������VQ�x+v��⮿��F?C� �nEm�Q[�g���l���)��s���^2��|O�R �4V���H��A�D=*�8rm���Ot8�``8M�y'adJZF�Iĉ�P:�v%�ib�6<�B�������l����>�Qa�6TКD����u ��A�)����Z�م���*WYh\�3����ʨ\��Y)��~c����t[�XZfsz�:*��M�2X��˦�Q����/[x�yA�<���B��ӕW��{n�3+������{�3:�$� d�Z�V�l�49_q����E�E�Vk憛���������k�-���i�
;h���a�����e�+����h����v4���|bL���G�ߠ�$�H�_ #�'(��^ү��+�����Qw.G�
��HA�; }m�1d�����M0�~�_���v��'�Y����s=	9�"���W��N�;�o���8������M}��|+��u8Ͻc v{P��Tﳇ�&�<�� p�"�#5�JGܿ.Nj#��Q�Q����qh��pw���H�= ����#�hD�������X������;q�/��`w�����C2#E�x���0
�|�x'�&���O�7�Z� ��8�uם����!����h���J��޸ǵ�ѽ��NW��h|�����k�b���%Uћ�Q9Q���6Yx���Ź`��7��=�	�	8�={N�;X���Lt�~��w�?��G�?O�c�8����Y-� W}
`��f@ˑ���BzA��G��i&|d�1��>M�RO���^�0��zf�OU��N2�dA��y�(���/�Ϩ8weQ"�5��U�u���=mv�SxQ�u��P3��[\��ql��k�k�P�"ڒ��0�J7��JJ�h�Q��G��l�<P(<N%���I�r�A�W)�cz�?��������U���YG��:��q�{��� �Y����
]��2H�z�u��I�����S�| ��E&ܲ���sm��JU�y�kv�3�=�r����ϳ�O?�Z|:��s9����"_�����ȝs�{8�qz�x���b:/6d,fPHŉf.��GN����=ډ݈���/�' �X]{qzHAv�X�����9���	�ð^�p�X�q3��z�)h�����q2�������gh����4�	��Sw'�F!S��.|E r��pV�S���Z�ֈ�A���(!�տ'�g��U9��m{"�uF�-1b	NrK�	Ă���۞�Ye-��A�=�j�6'�a(�(�Q" �x�������(���tD�5 OhĵZۀ�N�ʃ��(�CjG�@^�7���-hɉ(�H:7��OK��'��o�7�Y@ N��R������ęh�8��#��`~���.���gq����Ż���tf!O�9�h7ڕ>J噑s�n�Z�bU"��A�����1�#�#0���k`�q�?S�R�{��s��?ނ�G�+��$���I3���ǔ�@��
I����̓���s%��wk����y�9��*N��p�w/��\*�]�~��z�1"a�s�X�	��U\w(Q(�P�9���5�h"=(�r�C�Oi��#�����_�����I{_p�ڵ��Wdl~ͮ��z�k�^��_����q���a2�%��Wq�<\�<��X�Ἂ�4�� 2Q�+����S���'%w���d��0WD�v��I��,r+p0��~�3�P�[�k�r�lvx
v	nz7D�2됿��$��WD?��.rp��+>	���JE;3�eHB/���!X��Yñ�G#�K&C��d6�K{�$9���{u�(̝���`��^��]��N��_��O��l��/��;�ڿq����b./����!w��8E�C�	�%�� &p��pa5i�����%%e,J?��F��j�x�l�$��~�>~�Q0�K��'��?4���%��u�.��h���_я>�:p�<�y��Y+�.�m��bi�H�{X�Wg�q]���D�
��^�����F��ʵ� �L�nG@�#����'<G�+/�s�q"���a�������g�Awx��&U�r�p�}����/��,Ǚ	{���u�M�}$m��\G�ә�%�S&�S��ca�}rX�'?���Ҳ��Mb�A6qZ3�P�whF{b�x�gݧ��_�}���*��ИU����/I�����(q�?6f���ԏh�����QQ��M6{����W�¨'�Fm��z���
z�ˌčQ�����"�hg�E-4v��4�5,d��Ic��ٿ��nU+?h����'(��٭���7;+�O`���7;�ﾍT��;�d����};�c_m`u`�Ncu�΋�N���ٗ�s�/7�������v�?4�y;�w�]{�}��O�O�*��fW���G���>��_�Pc��+�_��W�����P��g�-d�ư˸��.i읷��;{��.j���Z壼՞�ٚ������Ô�5vNcg�3{Mc�j��fO��Nj��^��q�;�ǎ��ї+G5�������G�)G`Gb��a��^��j��)/j� .o����������?{�}��y���b�kl�����vk�]^�s�l�{v���lW�Ӈ�׎��-d;z�?jl�����m[�m�l�3vek {��~oe[4�4&yZc�=٦��&�m�`5��f���ae�ƞ�o=u�=�X^�6LY� [+��ؓ{�Ofk��(cM{�>���`�h��e����al�[��[��G��(�jl�{DcK5��O��p[���sآ�*�4��B�0�-��|/6Oc�56KcU�6�ʛU�R{E�����r�/����5�;��i��$C)��J��*%��++�؃�l��
�Y�m6�0��X��r5�3=H���tbW��l�M��T�M��L�b��g�$�L�c=<:ˏ���8��m���f���X���_��46Ə�jl4��X�a6�+����ϒ��*�lDb�2Bc�q7<�%�.�0K`	hH�φ��(�|ٰZ)6�"��y+�>,�V"����R�Y\-=��ء6%֋���Ÿj�(Cmlh-��͕�hl0X|���}]Y��B�sـ^m��X������X�Q�OT[��(����F�h����^mYT[�Zd ���V"��᭔�~�g�ħ��(�X8gw�ܣ{��Cc�ѳ{�&�(�4�Uc]4�ٛ���W�Y'o��oo%Dc=����'ł0s��:h�=t�^c�`�v����5��6��&���充�g�~vſ'�V��ʏ�b���| �O<�c������)���[ם��U�1/]w�Н��yBwd��ٸo��=4f�$V�YZ3���4����1ŏ1�ncs�H1��ړ;��4w�c���=/����WBj���>�k>�-˥E��\����u\y�Z�:]I����/%�R+{g��8E�%wD����5���!����j����wHG�1��l�����O�gGYN�d���1g)Y$�*����/�p�_XGv�R�9gK�����Sn���u�gp�9~4l�bzY�"i�4X�G�[�f�'�
�`+��'�e����L'[���F�\/+7���j��g
�\o;��KJ%�P��A&��~�>���Py6�N�H�M���-��G֘B�5�Ε�	���f���nr4��q�Q�]���R����B�|�wH�ѱj'o�����FG�Il(�̗���1�4CH)��K�|�1�n@O�1��6ho	'7)������R��9�tP�&���MLI��3����r�����y�1�� 5+Kq~�<u���_��T�ʧ�OXG��2��`����m0y��m��9�H:�͠[A�B8])�f"K�,�A�CN�栺�(�*�-�{q�r�v�P�[��U��ē�z�[��^�&�|U`���:��A��.�����o���R�>��Yղ�K�m�Y��F������ߵ�Ͽ�'�~LOՁ�d���k�tM��Ld_Э��n�ۻ����d
��۷�D'��@]���}��6����g��8��u�'ҷ4g��X�G�]e2�@T���.��,��Uzs�|K[Bq}Q�K?f��R��� �&ɔ��K����hG��4W�4� -݁�ס��Ć�{�l�0�B����O(�^_O{io~�Z��LN�{�tJ��m�Y|k�l5�6u�j�v$�B��:w���kLz�&�����}7��w"Y��D���Hs�%��1��C��l�<T�55���C��1����d*�*M�N��J�ҭ�V�UުlU�����Z�Z�z<O���Kϳ������Mϛ��<o}��9F�I��1��rL=f:f>f9f=��s�S���Te�:�4�<��'�9B���>�zG���SCC:�
�|쾽�}}�R�CE�lt�ic��ի{|��ǿ���o��yS��ZZ��)��vV;�]�Q��O��is�%�����>D��2�X�DN�z��α~�F�j�&Rc1��A��O�#F���K��ۇ�ދ�h{i�9گ��n�*�v��˻�� &9�mO��Fڇ)�ؖ�i��J���Y��2����*QkP�;���^�����hLx�|�_&��O����&zBH��c�ڷO����w�-Cg&/J����U�i@�ܤu�'�)��Z��cB�˻w�>M#�̫����a�{E_y���8�'�d%��?��J���V5��Ֆ��5j�j���5��M��uk݊0����� �g	�~��:0ﬃ{r�����Q4���ɰb��A`�x�A��fL3�-�?�����W��ܿ��ͫ�<�脣s_N�B��,��kO���Ν���᱇7�W\1�k�C���C�5��ʥ����L=�'a�3�0S�B�
�YI�YV�m�������x5_�5߁���P��	!ڑ�����`Ǿ��Z7�^�/_{�l�r�C�?���wh[h�1��5�]O�݁��M�֘|V����j�
�M��A,��	��b�F>e��k���S���õB��H3�q}�%�l8�c|�Ԯ}���ө�e?����޿��[{��}�e�v��x#�׾�����A�8@:��PSp`�5��n�����q������� ��3Ĥ�����x���V�G��w;��{�GP��8�<��:�I���4D��k�3�>����F�.y����꿥��o�z�oK֯_��ʁCa]����>���ݷ�-ZE����c�E�v�8���޻O��հg�T%}c�0�I,LV�xe
��4����)�)Dެs-^&�@����j����w$sC_���K�<�.�NRE�%�dXlX���tQk�z��"�vy.*�֩{�� oK����18
f�v��p�;�ݸ� ,�҈a&ctBK+WS*X��e+�=��[�ķ.~�Ē[5��5͹u���/�?w�t�fժM5�+7fv<�h�ŋ������s�>;��,�>硇��[�D��E�)I�ԉ��J%5��d�\m{�^�ִ��)���hp�%��9���Z,��T���+�X�<L�����;6��_n��R�u�`��pk������#*��M�g�zi�˔+anڑ�>H�7�E-�*�T[�U�\D�r��������=�vU�d�T�������cl���r�6Pl��!�v�P���Ŷ2co��+�Ij�Z�9 �>��[=���v�]Y���k�E�{�e/�2�DĶ|��o]�<_���X6�Mm[E�H/5�-�/�i�@�QaД�諢��\��կ��k��I�'�I:�v��}����N�:u:��ݺ�����Mݺ�58��ڛڅ��®+�ұ�ćt��Wk,+H��J�-&m�e
�G���z�s������c��1ԧ�������Y'��K��툶[���':�����J��^[���)�rRd���2|�[lk��Hk�?[�b�eB(�m�#�����z�2�i6�!Sz��\:V?�Ǧ����"l.g���t�meЖ�lV� �Ǫ��p'z��6L���~�S������[��VȠ؎�mIkֶ�}3{���~��վA\S�8y�hڥ������r>�};�i��>K������Ô=i��z���W��u�+�<�hZCK���{kt���wV�ܑ>�S�x2�B��P�Ц\?�ςL����s�z�۱�G7
��,��F֟��� �O�v�|t�)��6�H�z�>�],��k8�D�ץ����e��P2��b��,�7#����T�I��V�Ĉ�����$�XUU���$�Sw4��Gbu�B��g��ӵ{���R�@l'�l�����9�ҙvc���,�p$�g`��6�)_���n���}B�!��޽k�6i����,�x��ҥ�+���_�&�`�ɮ�9���ƛ��o��@�m��h߾�QWh�������[��\�y���6/燆�[?�#��N�i[�s�E�V���dm����
��.�W|����Gb{�$/���� �E2YÂ���A�2���ـ�yV�	�೩k��#���tn7Ы��i`HTW���]����JU�'~�Ś%J������L&�>@�7f���sER�u�~�nN~iʚ��O�|���c}�+�(ش�ꉢG����*�߸oв����z�/�����^r���e���G���W�	���1���^��t1X�1
?=�D�х�:E�Z�׵��ۗ������,�n�m��/N����Mv�"�;ȧ�D��-����
�_�6B*���[��rY#��mގ������m;70)~�����c��lc�������/pr�U_��W��sߐ�Ĉ�"�`�lH��H��i��OEY��4����J���bu���L� _Ԋ1��/���D�<o�
�p�?Ej�ii���s�Py>���$�;���a�6���jߎ��:Tw:�)��ȁ^VՖ��U�!��7�{D����S�n��4���[Hc;DG9�:F�l#��6i�u������l������cp���L(��}��p=�z�����m�K_z����O��@]7�����Y�O��z��,��C�R��̝����':<:�_��.]�ӣ�鲾Y�T?�ڞDŶ�YX�������vO_��6Um���EG�+�J}x��<�/y�8�u�<�7۰b٣�V=�lE�g�O����빛"jk��w�|p�҇W�9�Y��h��N��x���B�I����ض�՞��du�����^m9�7s_Q���ή�ܮ���]��&少�O��h��ߜ����>txϴ�q{���`@��W�b�^x���p���`ɮ�E!~m����͛��ҧY���p_�\/����³a;=r��n�$�X[�)���_��۬y�X�l��e�V��Ұ�=�1��G�� ��y�{��K�?���'z�?����oR��S[�j�'}%���Q�M���ni�����v��S<Z骺Ɲ�~�k�������4�t7���?;�7�xq��I�O������+��KS&�/�0�E(o mEm4V������m��C����"}�5;�����<��J�LĢ���~HO�:-ʵh���LǙ�����v䙹��b�h�D[T�]�=�{A��t���5�����ڽ���FȾƚ�%�Ԯ����n��RԺڛa�y��z�{�@�چ���G`��2����)}��/�c`K�n�'5�����q����&._���5+-���);3�o�Ԋ��ŧ���Tц�Zi�[���[����^�o��`D��}�S&�j�f3n�z|��k'�`�b���j�����߫d��E�H��kQ,�Au"�o��̊�[	��K3�dumm�]zN:�0R:X���jX��5옖�	��~̗��,8�G���)���*�Y�U�2�j��p����b$�IR�PJ�{����k����ZyZ}�5,^v����O�U�,��f=h;�*L�J�H���!���	�ȍ��d���й/�iѤ	�]���h���r���Z�-��#��!䏱]|�-��th���m�v�݉@���x�G��>��S��n�j�9j�-s�>��IY/����&���xgРk7ś`�oe�ã�(%J�2E��,Q�(�����04phۡ톶�ah�b�X^�,V��[[{�i��͚�5�kڮi����k�B�"H��n�j���x(�)��tWߤ��v�<��g;�M�c_�H��}�0[Z�U���7,���(�WyڴAC�}�h�;'��;���;���;�]�u�Y1i�Xs"�S�}I���_���?$@����������TP�vm�ck�>v��[_^�u�}|���|p��+[���Oq{���<[�����ə����ޱ�c�Q�M�$;�qy���n��wcxk��د��c�_z���|q.��\�Ö?�pV������}�-��x������g��.˳�>
��ѣޛڝ<�A�ñ�i�1�yr�!h����o��e�V�\�l�Զ禼�׿8���������2&���5ZӘ�k�}K�>��z�!c`�#>����	Gb��_:%N1`��y��Q�avb�vqP�O����Kb�0{�OI�i�4����6�Ky�}����-M�Տ͍�����w�i�^�I�m��/*��B�bcE��H�� �� 2q����V�����Î"�cک^�&�/$������v�{�	����[:nd�-o�=�\��7�l�X8�#W>V�v���3�d�{�{s��'����Sx "���Q#C��nY��ph�Ѿ}s&,�%y�[��;
Y�B�f���^�^�ٛ$>�����a���v_��`��A��G&X�|�k�|�|�]�2��O��ͷA��Ě�m�����4mb�N��)-��&+=a�k$��X������]�:WBc���d�e�z�^��n�.�� ����?mߕ���n�\�X,O#*ɋ톜H��6TR��I�������tzBQ~2��I�	��w��Mo����
��E�Q/~h23�,+R�$�sgo�MCs��D�tL+�
{L&���6������F}b=pF�Z����a[�1�M
�4�M�?��!�x�"13S�	���j1���a"����3��:�5�T?G���v������$�v�ڲ�r�������#�֙�T-uV���L��p�@��2Ph�mdK4'[�<F�ƙ�,�=&��B�/*3-y��y��K�GOok�̂A4�l�!�P�HC�A��	֙R�R`�/-bs�E�<e�u�5 z��ݎ�4ԃ�<����O�n�{a�>(p��p���i��߰Y�k���җl�M�l�����!Ylm�Q�6������N�����������3��ʓxY�M'}�N��{{�S���7�+�?�9�8����o�����`�/?;�������h�����{�O�O��O+?K�&	�J�����;�1<'$b�����O��9IS�𓴠��cLj��)������H�U�?��BBb}���������K��?Mr�xܲW�#��P�>8�)�Ljlw?Kk���U���S�i�i�	�M�ȞX�7V%�*��''$XшȄ��=r��uOHEj<����ȏyv�?��ۛ�,���v����ҺZ-���Y�Ⱦ���,9���[�L��'�v�/�43$��6*�[LX���D��ւ-�U#SZG���|��F�D{���΋߿��`�17N:7�7��x��%�ȗ�K��^���'�,��c���ɏ˵-@S(����U�j�U]8��)�T`���	�j�jg~������!�!k�u�u����<*=�yܶ%ت=%�A������޽�h��܃{p��=���܃{p��=���܃{p���T�'��=��'BZS���\�J\ߢB�wz]"2)m�v��v٭��0�*�"��:��ǌ��@�1Ꞗu�m��E���*[pwԚg�)qx�u��=�u��.���1ʨ���G�Q7��EF݃�x���{��l�u/R��a�es�gT:��tsDGE�vL��/���,��.w$��D8⊊�W�#=�"�|V^n�5!of��*GNAvɌ�
Gvy����QV5��0Ǒ[Z�]X�ꓑ]R�]ZR_Z�฼���GtD���s��?5z痖`�JL_PYY���YU�U�9y���3�"J�*#g>XYX��7'���,2�0'��"/I���p�%qt���sL�+*��-��x��Z���l�N�Qc֞���Z��u���,:*˳s��t�淤b���VŢwA^y�Q�]R����/�����pGe�#�d���������df�ӼgeA�a�윜��2t�*@�H״�k�PIH7�udWT��fc>h0��8��2���_Xw�� GFi~�l�<���<���4�*'O��-�`�ӫ*����J9EU���م��U�`��И��/�U	�U���	w�	��}+
����sF��;*�`�.���-��́lWt��:1����;p3�W��`�<10��QQ�>3/����:.�Kr�rJKr�1Vk&eO/��'$нH0��%��0C��ʭR���3GEA6���ghl�ɳ��YZ�(w����UlG�ܲ��lL�3��iq�\N��4�0��;ZvQ%\�������+�|Ue���r�*
g�6f�-+�����f�H�⧢�L����
�.r#Ђ�1��KE�XR4�Q���!Ry��"їW*�2�m\K$~��0��<��ҸC�ܮ��tC��`#:��&N�
v�B�*-ld,oN%V�#��K,{zQ���-S�]�(Ȯ ż��z�tM��B���
iWBt	ɲ�E|e�qCe;�x�zqu,��y0{�Z,)m��ݱ�M����9S#IcR3c�2�ǥ':�3i�c�%'$&8B�2p���9b��Lz�ǥfNp�IrĥNp�JNMw$f��'fd8Ƥ;�G��$'�-9uX�؄���x�K��HI��	��c�P�Trb'6:1}����'�$gNw$%g�r�I �H�K�L66%.ݑ66=mLF"h$�ljrjR:fI�!@hؘ�	���Gd�cP&���q	����G�s�@�t��.AÑ8�����O���LO���r�O3��hljB\f�TG|"D��OI�y�(�R�G�;�F�O�h��w3�iR0<151=.%ܑ��8,�W�����a��'tM�v��I�H�,��52"QL��o��L��
q9��1降��O�Hwĥ'gp��ǀ]nO��2��>��R~��x۝ށ^|�!`Bb\
fp6���J���WV�}�X�zx�T����k�  ^�����*�+K�<z�kZ\|K7�/�n�Fz�͝��(X�C	�G)&�+�J�6X\j�{�E��{!^faXE#���kC,+/Đ�兕&��*���3��rc�j)��%��yeة
g�͍@�r��	N
K�����TƸbh�c� ����E8�d��22���B2��J� ]I�k4��Fm:z8H<�T"��D�<�M�I8Z�I	�G���)8Hz#�
q��k���EO+I@m&(�#U葃�٠2C�t���;@��}��n!�90��f�g-�d*��h�*A�G)%�9���J�hpћ�o6�5�5�9�|ѪKTiH�%�1⫕s����?�Jq-?i�ǖ�"@#c"�l�� J�������e�Y��!m��'�$���ҍ�Fwڄ?�_ ��͕b�n�B�k�!~>�n3�z�F͝�;}�*���
|��~���-:��la�b���V
?�5^�di�^����:��,ϐk���D�c���/��5Φ[X��p�W��D�/3V�>���J��+tYrM�hV
.���l��=�C��.
���{Q3���
q�a�l��ǁ*ė���˧�`��XP�O\��G���㮍<6����kA�s>c�NxKp)f�|6q�+$��6O+�S�??C���r�Y����d���!*��6w�\�˛y��m��a��ux�X��e��[���?#Gx���"J9e}=��6��/K�Ҝ�mY�GW��&�f}��\�!_D�C�<�s�s��+��L����>�~\dDI��r�ܹ��B���:3�Q٠X*"C��cQ��|w�4VCE����Rv��>�!d�6,5�1n�|M׆ɳ���bGr�/׼��ڼ�\�o���vD3M��X�������W(ֲ+�q�+�����r������\��E�W�d�q.�r��^%nژ!~�����3�bh���w]s��Oů���r�yX����8�eN���R/w�1ܰ{�W�Q�܈@y���ft]-���Z7-w�<#��5��l!U�r�}1�Q�#x׮��m��Ii��L�ԍ�*c=�,1O�1��U{�]�w�lY�G��_���WL���q�0x�����Kw�ΟVY���B~1_	if��隭�ӵg7�:׊�DQcRn�hN�Lx��3���b��m��������RM7�H��/�7jjI�!�����]&�|2]<�?��@>��'�pǿ�=A�%N<��C�j�:�ȿ�?S�ǉ�7��'���v�{~7
�SA��M?��g�TǠ�?����,��s�T��-cq���	�F��R1*S�>��s����Y�s�,ftq6w�?�x'~�2EК �O��F>�Nㄎ8eNs8Jw�u,�i�g>nS�Ix�˒(8�-�s4L|��у�}���ϔi�ry�x>�(Ѫs6ư2�7Q�0t����?�q�!
�!��_��m�.�.�.(�n���B�8��1b�x�k��3��g��U�	}q�q��LqB#w��E��u�������RD��1Q�Ȅ�E��d!�0C�:M��u�Hq��0!#����5��8���R�+���$�n�8s�Y��S�k���ewje�X���W��uF����mp>���\vk��FΚ�׵�\�~K��i��nn��O)����u�z�Jľ�#�;����_��={l�J���p�k�3=
}�[�kj�㳾g5�y�s���\�S���7e���C�����=��y��V4f%��Qژ��O��t�4X,z���*ļ�dUƈ����2[d|���h�v��'�2�����J#3��U}y�������_��K�_���w��T�B�<��0����I'\�{a�-���}�Zi��r�p�<װ����Ӫ�=�x9�dr�߱�������m�e��H���Pi��	���fԟ����v鏨�v�����?Iϣ�Oڇ����P?$G��U�_�^C��t���|B��r���[�_�/�~Q~�w䫨��	���J$�k��	��H$[�g����[3�_+�G~$jBRJ&�]�=�D��-/"Cf��=HҊ�KdrQve	��ЄS�e�^�����f�����3��K��,�sr�h�3J��G�INu��>�1*�c��HI������)~��AS^9=W�2��9�"$T�IHiv���lM�Hg�kC�Z�W%���9ҍ����㠆+ݬ�[���gt-�>��N��-�B���Gqm��(2��������/#1�T 8�L��(��c��c
�X��%H~X^�+�ɋ��3���o�^�3�t�I-�|��ėt��#��E���UHO�<q�D91�����/��\�>i�G[va�Q�hh�霆[�/Бl�h�c�I��!�C�訥�BK��t�T|���z�~N���G�I�d��Rk��"u�"�>R�+%I)R��%M�r��R�4KZ =������s��S�#�j���)�tAzW�P�T�B�Z�)�f����|Y b�Xw���A,��`�,�Md�X>+b�l{�=�V��l�¶�]l/;����Uv����g�k�Kv��b��$�e/�On+;��r�-���	�H9M'O���r�\)σ����'��3�y��O>(�O�g�7�K�����\'+�(k��X��Zi��(]�����*IJ���d)S�\e�R��R(++�Ǖ��fe��S٣�Wj���)�rAyW�P�T�B�Z���V���6�WP��Njw5J�R��j���NT���j�Z��QRQW�k��u��KݫP���W�������G�5�K��zK�7I&����gjkr�:��MѦ�!��HS�i�i2l�%,���1�钴�ם��h����I��,���o5\ ��"�ٹ@�j޿��u�B
�6�xaW�C`���K3�e�E�9x�VP[!�M-��	�]�>�3u?mA#)�y��+_!�~*�j8��)�i���tk�\��!��Y�}"x��|>�z<�u�՞)�4�T`O�K�����p�/-�g����-1ǋ�i?,(�<��4�D�Q�-��-��=�<J�<�1����zg,�M�t���s �
����W
N&sL�h<Rd	�)�G��G�<rf	��hx�BKz�ў+��jj�7���Wo��_ߥ=ׅi���N�V��-�h۹�>����>�y����?��ڧ׵��'hՂs�ù&�"D^�
�|DhcAc�Ay�h�tV�����,֎M+j�N����/��h�S��bz����ꆗ�[�=pgiv�7�H���dڠ-��]�s4?>��Ӣ=EPp���9&7~߭~���X/h�(F�kx�_u��S���hҹU�븧��7ڟqV�>ӹ���9nx	x ���K1�Qh��_p�w�����Ѯiق�r�Ԙ���G�9a��_ر��9�D�i�f�'r?)��.��}��dox�?m�,7\�О�����\n)F[�Gi�!�9"��1'��!�)Z��8��#-<{��xT���<^�$k��@k�gI��`��b#������v��>2�oF�ؒl��<�d�{�xv!�yv��F�{��'_�';��˼�����[z��o��I��-O�n5�)*����-�|���?j�,Z����\ƂL}�����ʏ�ː���J�w���"���!D�Uɑ(�hǑ�ݝx�-2N�&d��'�ӧ�Uz��Mߧ�k�Kz�ޢ��$�%/�Oj+9��R�-��H	�H)M'M��KR�T)͓K�J�ғ�F��Uv�trP:"��9�M�tE�*}.�I�J?J����Yk֞���,��a1,�%��β���f�26�-`��q��mf��N���g��(;�α�]�!��}��f7�m�Ȫl�}� 9H�$w���~� 9^!�ʙ�Dy��/���x�#�*y��A�"o�w�{��!����|^~[~_�H�&)ߐo�����/�Oi�8��J��P�(	�H%M�LV�+J�R��S+�*�ʓ�F�e��[٧T�('�3ʛ�%�rU�\�S�U~T4UV��]m��WCԮj��G�Qc�$5EMW��)j�:S-Sg�ԇ����zu��Mݩ�Q����Q��zN����~�~�~�~��To��I5�]i���y��������\���M��X���]������#�,��HVF���w��
�d>�n�AM��n����4��2�#�?�BE�ԩ�x$W��]@�ɣ��	\�p��(?������UO	ny�eiop�R%��g�<H<�	T:"#��
�;��ci*�ne\�B��$�ǻ�e�
��'	#p���~��+�<Ii<Q��u������h�8E���@�G)�T� �t��e ��ZUc�� ��f�Zc�t��6��x��$K���S�G�h�������W>!�v�T-t���-Z�pGv�V���T���%p5�0�N����2��.LkE�.��Yg���Ch��}��lf��d��NQ���:�(�X��H{�=$\�{\��ϽK���TN��q�K�ncg��m^*�Z8�(�[$\>%�|�X�������+�4�i��K��i���i���2�u�3<&�(y�����<}_���S�2��l��	���5)�q��7��`<�X/��W?������/���P���^m�
�i�ĺ�)�x>êy�5@ϰ�<�a�C�r���O.���"��J��p����b%~(���z������Ur��?@Q�Ի8zJI���5J��3�Ūh��H?��G���=
��H�����0M�$��"�Ci�j�َʿS���XU?aY��3��� 5W�%�ޫ��ƣ� �3�A��]�ҹedD�W���%׆�����_3�-/e���c��R�Gѝ�`
�~K�$~��ƒ95AS���2��}i��%�Et��3o#�� OD3��� ����D�,�$�"���L��g�lClq�ؖ�L�w�dB��<� ��H�3�|�������Ɍ5f�Nl�C
���NRw)J�'��R��)M��I�R�T.͑��VIk��i��K�+��3J�J祷�����kҗ��T��bz1?֖9Xg΢� 6�%��,��c��tV�JX%���GY5{�mdϰl7���#�;��d��v�}��ط�G�ɲl��rk��"w�#�>r�+'�)r��%O�s�r�<z|X^!?.��7����y�\+�O����������M��BU�)�J��tR�+QJ?e���PR�Le�2M�W��re���JY�lP�(ە]�^�rH9����W�V�W>R�)_*7�[J�*�f�K�S۪���F��!j�:RMSǩ���j�Z�V�����j����Q}Fݡ�V���#�	����zI��^U?W��o�U�$��&�����)���a�c�1Ś�L)�tS�i�)�4�Tf��,�a�
����ͦm���=���Z�Q�)�9�ӻ�M���0}m�i�m&f�l3���A�N���(s?� s�y�9Ռh '�e�/pL��<Q#��K?)�ԭ�h1�����ϵ�>�{S��,w`��>�����\p��r��a}��n�MpQcB�����i+F����͢�o�[Eo�(w�~�:��=H�Z����}�h�������gq����O�Uw�C�����_��k�O�>�M��R���]?[�}��&=���cm���k��9���{���[]ؒ���󯶬�v��Wӝ+�?�z��ף��k�W�[Ư���_�0έE��!���3zn���w�c����;�(d���n҉<S��?�o�x���Ct��=G�O\���o��!$<gy��%��YE6���<K��nRKƓC��'��iRJ� ~GΑ��r�!�c�N���o�w�)r��@j�mRO6'U�j���ښ�!�Ӷ4�����P�"�L{��h?� y���~K�M�=qJ��K�z<��,�<��x�2�}������x\�LMy|L�����󍟴-�R���!R@����g��S���4ϴ�������i����n�>�A��	�ӛ�K�+����Mu�oM?�4�l��������sWs���9�kN2����Y�)�\�Ls�y�y��a�
B̏��7o6o3�4�1�7ך��O�ϙ/��5h�����k�M�m�����`	�t�t�DY�YY�-#,��LB,Q������̱<dyĲ
��Z�([P���Bًr ���b9�o����
|�������X%��������v�"õ"õ"õ"õ�׬�OsWT�q�w�{O̻�~�h�jԤ�PeǠ1��C���R��D��P�Xc���C��C�1���Z�d�c3��6Z�8�qk���Zc�1V{�ܧ^}<b��0��?�ݻ���sv���8�g�s���"Qwm.\��D`_^�X��E�!� ͈D+���ލ�}���#�㈎pg�/"�0&aY�����a�`�P����X�D"SΖs���\��2ډ��\F�ȫ�,� yb=b#b3b{`y����`O"B�Oȧ�3�y�<��H�D$@���0F�{1����G@=B!���L9���RX���B�� u[a;�;(�Pp �18	���E�� u���ԝ�*���R���_������nte��o&
�zJ>���QPsJ%�G�)�ԜRK���5J�Ҭ�(�3u��#v"Po
�MA�)�7��t :Ԝr��Gݩ�;{e����Tԝ��SQw*�NEݩc�	j���f��j�Z��U�U���u��R]�6�����Fu��M}_ݥ�Q?R�G��)��z^��1����%hIZ�6\��j㴉�m�6]��
�YZ�V�Uk����
m�V��՚��&m��]ۡ}���h��c�I�vV��]�%���궞�҇���)�=MOק�Yz����s�r�R�����Z�N_�7��z�ު����N}��O?�я�z�~N��_1�F���`6�#�Q�Xc��ad�F�Q`�s�F���Xn�4V�:c����ll3�7v{���C�Q�q�8c�7.���c�i�	f��l7G���8s�9ŜfN7��Bs�YfV���"s���\e֛k�&s����jn7w��{��a�y�<m�5/��-��k��m%Z��!�=V�5�J�ҭ�V��c�[E��ܪ�j���2�֪��X�V��b�ZmV����m�ZG��V��i��.ZW��u۵؃��{�=֞`gؙ��و\D��F��{m�^��FﵱW��m�_��F��{m�^��F��{�]�_��F﵏"p�g�B�A����Z��^�;���$9��pg���s&:S�i�t'�)tf9eN�S�,r�:+�UN���ir68����vg���9�v�9'���Y�sٕܾ���n��wb�{���q��tw�����n�;�-w+�w��̭u��5n��춸�n����tw��܃�����v��܋��`|8^�w�������o� ||qoV�Jܛ��fύ��Y�nˌ��'�����y;�����==���E�ɷDɫH^%���ͷ�r����^�)�S���=�ʏ���K/ʏU��,�oW[|�o�~��$�k��%���s�ⳁ^�{������ҺK���Ϟ{���҈Ϯz�~N�z^��wu�O��/�ƣ}����{�7}#���[)O�/��^�R��G�x,y,M����n㮣��M��hsD����]o��ש_���Z��F�Xy|�0�#_(|#����;Ū�g9�''*����$x@��7���G�����F��ˉ��y�g�_�zBkHWc�3]�I��(y�y�Z��6��n[�K/G�Zz>�ć�|X�m<Ny�z��و�s�xCT�<��WP���<���7��J��ы�_�����c�FH>�ʙO�'y:�I�z&c(��Yު$�.��#o#�F��.�����gM�Ϧ����"��9c�Ј/�*�gQ��B�ka��<�Q�f�7G���l0V�C| �����9$S9�tm��~���A�y6@<�x"�O���X��]�xWyܗVEIz�n��Ǩ��ttw%�
�)��3b���L��0�HbO@6�lⓈO"^@��x�
⫈����R���o'>��x�3�� ^J���r�|2�������kS}=v~�%b��������I>��l�ӛIyf/$^����x�1����xi���#��k����x)��(�}T�@*s ����z��'B�H#O�c&�!���a�X�����s�.��-d{�YVM��_a��U��y�$����?/)���I-9�8>VJ�&�")]��g�������S|^����*�B`5��h�+C�x�*�/t7>�l�Y����_��7�������o�=��W���WW�7�j���r�$�#��VZ-�L�[�?��y�2P���>�(j�Q��I�Z����M,���S\���u��_�*�!�Q�X%<�8�8��ļ0!�}&"���>E�����q��8��C�bGO��ׄ�1���8,V�9_$v� V ��z��q�$�!6��K�����^ZI�\��:�u�D�F�e��;}	�g���魭e}Y��{���.m�7h+�J�NV��G���$|���S b[̖�ZV�^�ȚYkem��h7���#�8�`��G��a�s����P>���c���3y6������x�/���J��7�u|=��xp����~�/46��{#�m9��b�ؗ �K~�\�����$�(�Q�%g�C2��Ů���,�x��G!�S�G����!���n�:Ư~*v�aOu�z-�����)]�Ko�������H��9�G�q�)��Aq�E�YNq�վh����H�e_����?�둚^�'g}��e,��>0}˞�X���Ĕ�B�(.4��B�(.tŅ�Q\�,�ͣ��<*+@�#]o�D�J"�3�
���g,��Ҋ��-`�%e����Y��3XViyi%�A��_6���\�s��,)e�"g%�@�⑧Gk���C��]k����)�_f	L����l���DbM�DJ����]��+֧�����؉��Q*�Wx�c�B�I�J"��X��\D��l ��ɔ;7�2�e�G�ہ�^�߱{�IR#�'{��oI���w�.L�uI҇҇aۗ����Sy��;"en�=@?�$ض�O�k"�d��xx �I�<��7�[�8|f�L���̃'���x�������<�����Uxބ��m�3���_�����	w@0 ����w�0���=��W���E�ܩW���Eb��]0�������|XO��G�c�)���������p�#."�M�����/�!4������n�\��A������`	�a)� ND,0-X��p��XB�5KiGdB6�@@�CTA,�%�V�J��zh�Fh��06ɗ�sr�|Z� ��0�L�
$B�X[�B��,I�Z�1�1	"�����������Tf�V<� l�t<�bz��3�љ-t�]:s��D�(�����Q�٨�����}�;�[���g@��K��V̞�߻�y{�o��8�i�0�;���O,�
endstream
endobj
20 0 obj
<<
/Filter /FlateDecode
/Length 446
>>
stream
H�\��n�0�_�\ҋ*q�W$��������F*Nd�o���b�	���93#�v���a��O����4�>��x���;�DE���Y����NTD�p������6*���uwZ����=Q�;�.�L���!��m������J�k��)���~�GE�}\��sd����O���E�1��:���?;ڔ�i�ī&��o�Z;���mH�e�ܪ2��P/P[�5T��@��PoP8Sb�PP�"4Te� @�� `B�P \K % ���A�c�0�+�aJ�
��( S����BKj�+P;Z5<��<�V<��e��E8E7ܮܮ��]#�]@�Fs�&�|&���f�<��C��i5,T�a�4<�-yh+xh�c�a�аdhX��Vd��Wg�i(��e����B�c�F=��2i�w��i�*}�	0 �k�
endstream
endobj
25 0 obj
<<
/Filter /FlateDecode
/Length 14523
/Length1 34888
/Type /Stream
>>
stream
x��}|Tյ��g�s&���+�+��1	I ���$3y@�g^��O�(-�"���H_������U��j�����R��ZJ�3��sf2	���~�{����u�Y{��Z{�מ�0��	�2WQQռ�3��`lS&�fy�Ug0V_���Y�e�?~��q�+fU.���(�a�n
zY�؜;2���1���6������|������]��z���Q�݉67��뛯?ecig���zw��H�~2����u3�X�1��bL����Ę���K�Ml "�0��=���ܺ槏��n������W뾶�5�0��.�?ov��'�j�~�Z��ޫ�8~�^�m��lmd�c�T������?�ؠ=��ԕrő���cW&L�������O�����oko�T��UI�s4�A���f�����Q	c�f#$�$@"�%
�!��EC}Uy�A�8퇸M��ⷬN�NG��UEQ?e�����B#�cy]����+ғ�d����?Z����������*3��}�����l��_�'��,���c�3�*v5{��zVǶ��-l#��gx�U���LG��l;���c�Y�X3���l5[�v#߄^K�
6����A�T�����l�.A����� �}�5�[��c��r��Ħ��!�5{��wa�'X0����լZ����(����X�}|
�ɞace:�;���t�NL�N�Cg!��b��u�3ţ_��;�H�)���V�ɦa�+"�F�ηB��v�m��o=�3������قv�> Ũz����9���5�\ ɰ 0�����y	�&�W@��e��@^�=���1�u��@f���>�=mcn)�zքՙk6�|���Q�H�\��m �ɒ��&�MF�ޒ�e	�hd?bqH-�⠼ne�a=&+$���H���42Kڰ�~0�!��Eb�J=�,�o��Ϟ5�#2
�K�WR�+��Q�ڜz��V��"�m�tɤ�K0>�������QH]��z���4�A�&��XV�R��X�����Įa;��> �
v'r5���M)��-�B��XqO��MH,��+f��4��fX�\�S�/��^��N���&ȿ�5�?���H� � ��[�|6��G�)<�M�<#�� %���4?��>i6�;`_(�|e>��=HT��7�hWr��4_��p>�s��Nl��=/�ڐ�c0b		�q�����_ �>��"��[�������i|9�TƲd��y+j�*q��
q&�J��Tc>�9�΢�>���������y(r��ٮ�+�!x�f�7&�Ƽ�\k>Z`&���������y 8Xz]��3]k�A�?�a	�c`Y? �xV���l��K��;�V��k�K�\�y,���f�,W��A�e~���͡,s��y"[\���ja1�y��@�~/��Ʒ�������J�z=�K�Ǟ��%������C�@�(�Fj�n�0"�v�8���yY)R2Z_<c���<�x�]����r̃�c��$w{`�e�E7����� ��M�4�ڒ���#m�7�AЙ��c�܇�f,Jt큑�c,����]�m{��)2��x^)q�Iʕ�e�����}Q�N�.�؆��~�� ���$?$�z��R��06mi������Fy�2�A��,s�\`�ag�6�1�+����8�����'�M�3!�c�<V-�a_��+ka6�[�վcԃ��܁�.���A����|��6И�>5l���b�LC� �_��d������ 3�&�x���|�>��4=4����H���lv�Dh��w����l�(f��y6�(�L>��"M��x�5�Q�i��G�V��?*Y�V�1��h��@7��y��'�Om�>g���l�i%��#U!�OD~ũ�eȃ@yج@Zپ��a���<6t2�W�U����I(5@[�?tH���ex�[��O�/1�5��X�R�Z�Ԍ�y�+g���^�0��v$�h4;�N�t���F��@���eρ����H�l�W��4)>7����@�9uS�<�j����SaeKPW=�����n8�y8"�L�5��N�y:���� ���Y��Y�!]�%�%�9Uu�ё�a�HQ����U�Y+�
�n�|KE$G�T2�:%/HYFSQ�����ETS0GS�z�|e���,��p����K��=:6��*:��OEg+����n)!�^ǎ�;ͫ�	��P:|���q~�5�Jj�������R���#n�}���m�;2;Ts�9V/���^��'�/t:r�您�&�u�����8�5�%�W������8�\��F�>��}����w╸y��K�%r���V�E��4vg��6�=����?O�G�%L�y_�͵��ﳿ���~í̑���:��`]cXL��f�ف�cp���cNFl��+���y-��Tc"e�d�����&�N���l������+�%|{gF�?|/�H�0��3��X��*v�4(E*F�:�}C�H\ӱ��e<D\��7h��������#�t�9Ң�����ܟ��V?^�6�6E�=9��9���C�#pF��>;&�<0t�!��ᚌ�Ì�����G�Ɗ���#�𝕦��a���b���'Q-?c�����aDJ�]�R^��AZUcv�A�Y89:�C_��ڕ*��<;�jHu?�L�8<H�6<+��Ю�]������Kdz԰g�~�N[��7qz��?�]��ߐu���ԽE���ڳ{�����2����I9���R�� �W��`��!��oJS0�yB���
e%�����`�:;��6:���{�S��_	Nt�n�о�%o��1����w��2��L��x�>��qj���t���,���8�A�&b���ǚ��%��6��T~	�`�?S��}��eI�]�D�;����tւ�礒�_���}UR	���js��p
���R���I��5|Mx���MJ���8n dk�t�|�4Z�6tR-���ɧ~��;$\)�뎋\�	G��Tu>�O
�NeJ]�[����26}I�Ys�b�٩H/���f	�n'�{'�G��}n�.C��Ɍ���وa7��fx�X�JG�r��n�"<j0���V�#�������~���:;�5U�~�}bڌg�����ɨ]��i&|�g�;�o��g�z��m`���:q��� "����6&��,P���@
�2g�1X�Y�+�����e':lCD7���81��^5R�~d���N��T�9g�K�e��1��Ӏَ�6o�9.�O���aׂ�lH;���>-G@��/#@ehN�l�J�n�P�]n�CgC�I
�� V��Κ�S��)D����V���|��uX���R�� v�K�$u�����!��^�B�����R��c��VN���FB��� �H0�t��ѿ?D��0� '�r2$�����`m|$� G�!٢�NJ�)įa���r�.��_�/a�#.qw[�	-����Y!�w���@�AXQu؋�,���k�8��~�z����?��M�ʍ��	�V�6`���wC'��5�-T&W�}�|�BW�r�S�Y�����k�Ѓ���N�ޑ�Y�a��l�?V~F'@܍�1&�Ӑq�Ǚ�����~�����?��!�;�t���z�w�0����ɷ}5?2
�O����X�л��lV%��׈^��k,��e��m��B��ۼJ��~!�pX�ЪPS�O��1+u~���V����U����{�!N���]��p�](9�c��K8�ݰ��$��~�89�?gQҐ2=C���Q�i ,�xa�U�l(���>� >���ceXUW"��B�O�g |	�a|�s�9O��C�M�����f�ng�u&2=�`����G!ۙ� 	�!�E.�3���U����3E,;���`/:)9��N��\�E����쩱��!�*����D{�O#$դ��ˏ�f]������g]S��Y�+�2��s(w~��Ń�dv�u%:\�X��k]GB��j�����6��sH6�o��`L���jס�l������F����@�Ѡ��a�W������u[�mC�ޖ�:�Q6�5œO�'�??+~vV~|�v�I��,�X�xt�x$G<�������Z)�z�M��_{h�ϊ�!�=�Y�g�}O��]�=�Y<�A���m�b�7W�I��c��s����{gi���#�WsC�?���%~�'v�(G۵R�(G�4�=gŎ�⇦��S��0�-U�e�����)�4�o��e����d�q��D��d�9Q|�.M�^����nzR���nY�mzRlڠ�r�0�e�\��a�����������zsĆ�zi<�^��mb�G\S)�ūs�:4X�#֦�5@��զXe��`-�C�����*K�Q�_/|����I���M˴�'E���q�ִL4�+W��Y�h�������{DF�K�D�1E�)jL�^/���
�Xzy����'�%9b���Q�"���"S,�LQU�ԪE�ST�O�*������Q�(�LQ:ϣ�n�<��sM1���6g�(�%f��Ί������V�^�3SE^��,G�H�N��.5��iNmz���S��ѦnS&;�)}Ĕ�d����N���M�$&����b��Tm�\1~\�6>U�K9��j9q	�/I�cSsS��16Ud��&�d&icz�1G���X5st���$2�(w�G�k���#�i܍��Q�b��!w�:r�� ��CS���b.�抡P��T1$Y�H��s�`�xm���5^꟬�'�pI3�@4�#$���zi�q����뛤��%�Y<��I��&����"55Y��+R@.e��=I$O�x����#�s���"��9"!�ZKX/�q_-z�L�4a84#M8D�1C�I1��H�0��$�Uu-V��~��>�j�B;�Yn_U�&��Ci���O���G�������6��3���C�A~;;�]�J�x)[ʮ�C�p��1l�j�!8#,�[-e�վ�)ԍC�\�:�jkT���D5����������e�򒲅ak�	MA�u��^���B�t��9>1�.D�C�)�����V#^���0Z�a����uT��{�}�^g��7��l7���*�b#�ѓC ���eyO�g�*�%b'�͎�u��9u�LW��)e�r���}�.����z2ƻ����WQ{���$���a��mn8$�/&h�[	|ǰ׵7�KqV��b�(�������z<�N;��A��4N
k0���Ā�/�P�2�(��j��=v��%,����'�{%N68ip��ڃ����m��3_�����/>�,N�{b���1��_<�"h���bN6J������7�єWm}�N�}YVn���/�/zl4|�����k����%���!�>>}����S_��χ�XR"���')�IWz'��3q�:�h��5�Y>�g-�YP��d�O~���C��;����1t�y�(�u����"Ҫ�bj�aIlDno��pb��Ǵ�=�XBlzO0�~2i
>�����a̤Č!|�dg$���}�A�V>��|��<������q���q��f�4�"k��+ �@V�;�q��������|���-1�4�KR�R;����ڏEa?��sJҔ�ܞ��Ab��E�	<AI	���/�IC&N:GSz�Ԕh�5q�Km�{�1~��`Ɍ����{��
x<x���x.��Ia�͟���0C3ۓH_��
F}9ِ�$�������&İ8#�����c9����'s�)�����-�~���U��}���U�4���^�K�5�2%A���F0����$��pe����ǚ��o!�]�~{!716���S�↱=���i�u�9�b�8���?�9tvnR�"�zWx���a���گ����_-NdK,��r+bb�+���ʥ�e1��ޢlPr<��/��3���c�$��'���M|�Ml��n����X�sO����s �a�q8��~�ز��⪪��ai�Ԇɓ�ܟN�$���!��G�5�?�kb]�l9;Z=�Tn�{��R�Rl���`Fz�~�pBK�@j���ib�1<U*����S����b�/�yXF�bJ�UW:��\p�ǚ5����_�6O�%�=�4~�d�17�כk�&��F�<g��)��>������Ĥ�Z�^p]�z�ƥm����1��ï����+�M�14�ϠĔ�"}Db�1p�1\��εO�%�&�W(ڗ��<�O?t\��{'��i�w�:8=cxR���g������Q���+�-_������1��߰�?��ה�([<��7���2O�,ZX>c�%�������	��%U��gz��-����,�+~��M�O.ұd�#m����o�7��_�iҙ���j��3�qv=��2�E�x�y���Wa׿;z��MK��i�� 61w ��%�~��1��[y�裲%')�9r������D���9�����S&%b����K%P��Ç�������}~�sWӕW��\ye�xF���ɽ�>���<{����ȑ���xp�U�`�ldnr|���cɢ!�V�θ�)���8I����ǒ,F��8�yo��Ns�^��q޲�e��2Ǉ�~d���x1:33oFFSKG�����Ɓ���I�t���$�^�T��s���i��ʳ�Mo��z�t��t1]L��t1]L��t1]L��t1]L��t1]L��t1]L��ԙ䳞���+Y�/19KĝUV���vY���U֘�Z��z�v����e��l �c�{���޲��l<����j,�ƭ�˜��#��b�s�`�"x5���Tg�]�Y�3L'��;�o��l��Q�ܣW���.ǳ�3}������V׈ڑ����q�������`k��n�t��f��\�*����U^OV\�w�{a�����R��������o�ij�uy|��Ɩp�JwK�5���s���<��`��ŕ�5n�Հ�zU�}�|-�L4������~U[V�������ެo��Ս+�6�x�k����%��ޖ��H�&�H��<�A��U�m����d��uv�n�E9���1�����vu�,�Zn���X���u�W�47�vѺ��b��������t� <�A`h/���s�[ֺ��t�մB�Ɩz�R��ek�מwm��ُ�Ԡ�ԛ,M�F�K���1���j��mk����[����&�xQ�\������y�H�I���<m�^I���k�Z���.21K�Mm�duck����47�Q���J�m�=���j�J���2��Ȥ1�����֍`�������Iѭ���@�|��v�i�k�`@���񹂾LW��f����0���`�$P����Hr���U��]�[�XV$�A�����4+�N��\�7����Z0rw9}-������WlW�Z��΍��,���6���f��������
�CD����R�/w |�5�r �7�X�"٨oZ�oR'�Pw-��G��`��,��X
s7E�F��楓"XliZ�j�b�)�w~ɶT�2in�K���Z��<AWzd-����
W:-�t�6̎��VQm�<��|�ƼkZ�j\n�K�]��
K~P�61�VW�;�ޖ�z�p��q��EZ|�w�+閄�� �2V��:�(���<�K���]��]�������V����������]�**+�rU�U-ʫ(tW��+����*q���ZT\5�lA�-*�J��ʊ\y��]s�K2]��������
W���B��Kg�,((.���G�Ҳ*WI��*�*�]mRŅ�Dl^a��ٸ��/.)�Z��**�*%�E ��*ϫ�*���$��U������4
@�������+� 4��|qE��U��Td���"��p^^��L�"W�d�,p	�Թrv^I�+������0o�%��*-�G:ZPZ�WU\V��/�(y�%�oefI^�LWA޼�Y����P3[�NuP�Y���y%�����T��+
gVɖ�=4Q"ٝYVZY8h2�P��o��L�_
q�NUYEU��Eŕ������Jb�����|�ɸ ���+���9"ܹցV����0�+��s�º
��z��d���ܣt���̔Vk9��,\'��g�,��X�sqі�i�_r�n�F������ɕ`}�ș�nʕ�m��g�{AwC�H+�Kw�#lv]P��hD�Ձ�V8���@�:{+�[Uw	h����A?v��Uަ�Yh��Lr�؂(��]���uj؇���%qG���c3�A�Z`���5 xv�����5�e#�C�-\,mZY9���E3�����B)O��8���
�;/�^�Y�A�8V��
PX��ТmݠR/[�P&�.Pi��W�4�w�یTםN��B�U2��C_ZA��I�9�c�ԅB����H����zK�V[$m+x�*����n�
��·k �{e߀�4K�D��W����c�T�wj����DJyYQ��a=����������4���M}m�����9Ȓ/h:�Ȗ��(E�|�����,��&�]�"s��E��w�Ym�Z]	�v�m��d�^���i��Y�媗��H{�H:u��͚a��2%_>�a���ׇ5�T[�n�Va�Rkk:L�Ur�uE�ѪVZ�ߦ�@�-ޛ��4�Vz���˙s˵@נ�}ܶ|���*�%�VY���ɶ�;G OA��b-XvN#v�0~@Fi�|vr��J[�G�����<B���j�Y��b�d����!Zm�4K\�Da��.Viq�&u�5;Tn������D��o�#3"�X�\���,ڍ�V�����k������nV�)�j����4Bx5�I�bK��#!��)�m�^H�im�M���P��#9n�9�*Wg�݋^�擞�s�}Q����ϴګ!إmx���������n{�j"~;lk�6,O��|����Y^���٦6k%�u��.��P_�����r�5ʵ�h�{���,�ũ[���sΣ�.��(���@�-��%�HNi�Z��Q/_�G�p02R؇���X���~��*S���t�0����qpaN���]/��1Ӟ�&ٯ�^=`{ �䯹�0&���龋xm��2��T�?�<�bzD��=�}x�M��6k�t�gj��E��f���L�Bm�y4F1Y���Pk?�����g�FzDϿ��WL���.y�<z�E}��XҝχSm�EF�+���Jz�9�G�lЎ�]�$�U^QA4Eb��ݣ+E��蕀���Y���w�?�_x�o���^#���X��T��)c���q�pW�!���u���|�u�^����%O�P}�\��P&�e��.�F �^�v�{������E}Y��P�T�ZVH��-���nG=�UHpO�Y��Qk�R���l?O�bqZ|�]�*�#�9���
Пm��v��G�gJMQ�4�g��i��Q&�3�Q��#�\��KJ
m>
lnK�E��d)�X3aq4�r�M-fѫa$4R��2SJH���4�\��8+�g�ʝT�l]Z|��+�#6@��K]R�*`����~�n�vfI
�"v�@ʗ'�P&Gȗu�E�gI�eEԬ̔��y#��HyR#��$L����:�#̒�JM��֕�c!�G0�=KYgں�hZvo�DI�vgJif�c�Bۦ��Ja��S
k�l83Jg��_j����\�I+;W+��Z,����\WF�P$��<��Q���}�E8���:
��.�â��H{*�9��h���Z���Z�<�X����;wt���Fǟ����FG��%�6wk׉����gu�y�c���\�S��wF��������(:���8݊�����?|��d����ӭ�`�l}��q-����iY�[F4Z�<ڼ�������5�jYn�#���nK�u�NŁn��o���,ߦ���o?��T�R�Of�t,|>��	i��.��۬wZQ�ʺǡ���(�=��[߫јq���	]+ߖ~�7W),�)���֬x��wz),�	�ƕM�Qڡ�@��G(�R�f\�F��	u���(������k(���@�燌;?r~���C�G�b���3FR��*3�d�3�����e���]�6��f��+Yy���bK�ܭ-P�*�	ɿv�J��+�8�++���q{�s�
�b�+�����H8���T���y6�rn%A��C�5Y?	3$�j^ټ�Z`|��}Y
����_ϱ�e�l ��Ϧ�]����l�ڂ�t=,G��;����}�n)�ei����S��� ���)-WVt��иz��e��(g�4�l�&N�;���$�׫7�*����҆�.���Q+u>�2u�,7��� gςR�	'B�%�#z�=�8�푋�c̚�c��B�Bm�̕��=�5��Mnǆ&9�������(\y1D�,KdR�kՍ��9�s[W(���e��o���C�?�O�
St�Pz*�J�2T�d+��J�2[)U��%�r�NiR��Z�F�6�Ne��S٭�S*�)O(O+�T^T^S�R�S>V>W�P�Vڅ"bD�H��Kd�L�#&��@��b�X*jD�h�b�� n��V�]�{�~qHO�g��eq\�#N�O�I�8#LUU��D5E���#�,u�:U�U���B�V�P=�
կ�ª�k��nu�z��W=�>�Q����_c�����~�~��RO�g5�隡��R�4m�6J��&jӵ|m�V�UiK��Z�֤�5ڵڍ�mڝ�6m��[ۧ�ӞО�~���������}�}�}�}�������z?ݥg�z�>Y���s�r}��T����U_�o�o�7�[���.}��_?�֟ҟ�_�_֏���'�O���W��t��8G�#�1�����r�wLu�:�%�
G��
�Ǳ��w�r\�9*t��֐�k� 6H[]j�ڕ�j��К��T<��^���fu����%`��Xn�R�9@�G�omC�������3�A(�	�F�2`�5���PPr�'�0/T;�G��j�V��#1�3T�';������
����fW��CtB��r�R���ArM������e�:q�A>��^G�בE��� �v$�Q�d-��RI�D��C� .	�e�K�Hb�$�Z��p��,#ȏ�0k��P.�iY�� ?��IB_#a+� ���W��@/eM�N��W"�;�Ur����Q�ud��Av��c�Č��L�|P� �|&��)9�P�A(��C#��B�0�G:˰+�L�E���J	O2'`c��v<8Ŝ����2�{���q�Z	�5�i�%,6�4a��'T��({]I�d{�|A��"mLB��y`�m4�/}��P}7���j�ar���煯v���D|���L�J�}���,	oo���6�-�n�����n0Orn�/��_�&��:^�@w��t���<�H��X)�\����Y,�ż�?����=*���?�--�� ד,�|s 7ǒ��7XF�J��_Ce?�4&W��$������6ˤ6>���I������W�B����x0��Zhu�F�zFYlN�����I
�IY,�S��>�/���s���J
~��q�"uB��e�/�,1���3��g�42YИnLg����=��7N�O�SƟة�ʾoG6/_0�٩St�cA7�Ga7L��l7̬���0�k��c:#�X���e�v�z�z�zbu�k^z�,���޽J�N9�Yo��߄��_YH��.�["ĺ�zK���mV��4�����TLx:�?�_�y��(1J����S\J����(��J�2G)W*K��AiQZ�u��fe��Uٮ�R�(��C�a�)�Y��e��rB�D9�|��QL��8�(R� �.F�,1^L��H��
Q-��B��*q��^lw���q��+�G�qT���7Ż�C�8%N��*Su�P{��j�:T�f���j�:[-U��%�r�NmR�X΍�m��6u��[ݧTS�P�V���������~�~�~�~��k���k�Z?ͥeh�Z�6Y��hs�rm��T����U[�m�n�6k[���.m��_;�֞Ҟ�^�^֎k�h'�O���W���U=NO�S�z�>B����S�\�H/�+�j�
ݣ����*��z}�~�~��C�W߫�я�G�c���W�7�w����S�i���9t����Hu�9�:F9����َRG�c�c�����8�8�u���q�c���GX�1�#�ӾGe^��hW���BQ	���D�T�}��f�UWF�k��*+�4�V�A��>G�8��f���:�<[����#R⇵^��F��I@î��:�?����"�QT�_#���e�4J�J-ϪC ?���S�G(�b��I2C�lQ���T�k}�k�EFO���D�<�F1��e�`�����M�JX/�p���.��
����<�e�é�w�B���i�kt��Ҩe���<��3�2M�5�p'?>^;8Y{p����x�ܥ�����f軥�p����7��U?|����(9����M����*E2�T�"�c� ���L�O�cy�|��R���_�&Y��=����Ð/���g��K�i���Z����|�� lRjh�(��P�{���'��P�D�0M#���`��C�e�VGZ�h��tj�KT�Q�'�jɥd	�7��(�����t�v�Q�8���IB����(����H��Oi�Ε���NU�Wi��,��/m<����$�%|_�G���r�}����$]�'��r����)��5I�E�Y� �G(���	q�Z���$�(a�N}��ֲq{�����3�P��DW��x�J��sZ�������z�N��Չ��I�l?�n����O+�q��G��'�Yr���VG����(�'~��"�ڥr�x��5/ْN�\�#0%E C4����yP�'�dI���Q�u����g��veA����P�A���"ye���u�Ͻ*���`� ˩�~鰤pVM:W^�Ԩ�BΔ�_zԇ¾TIц��g�����t�����!�����|F��/R_D��#�őj���&��*A��j�q���������q��2���"�P_!/��@�q-3���x"O���5�g��|*��E��W�j~����W�k��|����w�{�^~�?���5�����_��η�,Ҷ߈�G%�(�:	wI�#�M�9�skυ�C���W����<U��*G��!aN4�����~]4Wߥ,)��.�M�f$~������|�wI�>�O�$��e1\����)�zY���PQ<�q��C@���b5Q��b���<Y(GN�kO ����w.��d.Nl�l����M�4����o��gF�@/ley2��&�|�Ϧ��T��_寲���	��ɿb3����r�Y~��+8#��8sgV(|�ϊ�Zq+w���W�'v�z�f�f������V8�:�f+oc-�}�}����|���?u��������1������M�����ZzS�|���s�����-E�A��-iAnE^���f���[��
�y�~�Cȇ��B~���I��!N����v��>Ȋ�=?�����z����ٶB�]�i?�9Y��/���v�}�Nb�9���~��Vq@���_�oj���*����S#��4�y�����࿩=օ�+�>��$�n)�����8C\���c�r�����D�4�m�3��Ɉ���L��T���J��%<t~hq`�q�{�0���/��1G>k,��������)�a��F�~��O��>s���t��"朙W�b兕倳�J ��j��Z>���O k��j��F>���O �#O:y�#Ùy:[�z�dOSc=�Q���f�-��lnV��mb%\���4�� �l`���~fi�#�-uI����	��>ϴ�Ͷ�%�';u}Ǻ�%�Jq·�g����V?���u�)����8�8?���(����q�#��7
�"c�Qb��Bc�q�Qc��
��h1�*c�q�q�q�q�q����f�0v����~�q�y������ί���8C7⍞F���4�~F�1�e����W��35�=�����4��H=ܘm�UF���Xnx��j�1�167���Ɲ���vc�q����g�09۝���9O:�8�0#�H4�f0\F�n�ŨK3�
�
X�r���8�(���)��^���O�~�|�2���"�r�J���Ac�q�q�q�q��=c�q��/�=Ə������Cο;������_�2���H0z9CFc�1����Y���d� �gL1�����`���CP����ϒ��QS`<
�k<8#RsX�<&k�5�T�I˕߄���2�G�%�b�Q2�0�4��q X-��<l[1>/^�������#�����ô�
endstream
endobj
28 0 obj
<<
/Filter /FlateDecode
/Length 263
>>
stream
H�\��j�0�_E��P�:�F!JF!�}�l��JfXl�8���l+t0�-~��B�Y�=wF`�����(��]�Dp����a���Y8`Q�oK��3�����K���� ��+��Lp�j������h��i@���*f�e�NŸ�1j�2>7��3��6���	�^�	�>��@}��4�_�B�a��§l��$S��'���JDN�]�nD�,89�YQ͂��,)����>R�i��%���8�y<��޿�Y�T��
0 ���q
endstream
endobj
29 0 obj
<<
/Filter /FlateDecode
/Length 804
>>
stream
H��WKo�0��W�\��HQ/��e�a���+�aX��?��WV�n�8�hY�ȏ~�N��')$TߟPr��1<�$�A%��h��XV�B��g��Q�񭙥����c���w���7����8T���!��a�5�1�C�0`��i���x�Lȃ�{S��^��x��xxĲ�i���7�y�n�5܏���ld�P�K�lҘ�»p��QPB�lFj>=�@#)�ړ�9�5��/�b��ڃ��)���u�<��/?�:~Zms�/����Ez՞����� ��_ȀAN�5r�c�韄̯\j��v�r�%*�h��UB�B�zq߅/D��)�����=`���B�tQ�)�����B�|�2�+�0�X,t���]�� P���G� �Y%�E#�߉���t[α�S�<M����jŕÕ�X���}�Q�dk��,�G!p&g�`��`5����颼�UqKxB�KD/�SZ9W�Ĳ�+�%���)�4�����o4N��H�dYt��5�q��'1�+� �Y]
�UBn�,�4�k����E\0!���=r��G(����;u��v(o]E5���=�!J�2�yp���+(�Z|�
��������~Km�� ��ϰ,m�����R�
��2.4����n M� ~��Z.�K�;�j��O�&�-\�EwE�-�xr�]l�6%y:��r}�0�>'�!Z�r���9d�����|�������
�U�K��@^>5�l��Y���|��F�u}��h�Q��l�^�� ����!>��5̝��?<]��+� ټߣ
endstream
endobj
30 0 obj
<<
/Filter /FlateDecode
/Length 620
>>
stream
H��Mk�0���>2����mr��[)=�R����:#y��v���Jf���J��˯q�y?y���l(h��֏�~����2!x�C�C��H�������o�����2=�|�Z��Oj������'yΗ� /m�4;�4B�r��h(�W��]YD�0��XW�̶�yɊ�d��3Bޝ��K	-[��Y�����mW�,;D���,/ǥ42�^A�B��ɑ��@�����Df��&c.;A���li&����I�wE�[��\_�I3�G��6mwAf:AD��1Y/B���W�� j���X	hWyW�»�#�/K���?��&��_rMA�:�:�"����˝��بۖ�H�['�)eH9�e|� {�i�w)#g!���CӋ���LMe��.X��������e�5�U�Vl=�$��#YzQ�J�����nT+8�����]E��{Eвՠ,՝�W���&VA5̫���O΃�F���M�o�z� ����xl�s]�<������$�-��9� �8t>+CIiI��=�yjP+��K�(og�݋�d� A�{�noX�� mA�~�s��o	��*]z�{�Q��9�eQ�\�� �	0 i��
endstream
endobj
31 0 obj
<<
/Filter /FlateDecode
/Length 676
>>
stream
H��W���0��+r.��eٖ�t��Co��-=�R:���*�i��nKmo	!�쉟��'��[��N��6+�8Îp�x{�<ޖ�E��V���f���bV�~|Y��!���"ZM0*M�}	�����0Ni��[_����η�-��M�1V�z�ʯ���(�=ݾu $��A��0[�� �2cG�$lƒMbǵp��o���r]��8�y�!�j��Cu��!� K�qc�Ho��e��Ρ�h��_וc�=��(�
�l��̱�S�Ę��<r�(�|_x �Njf��Sйj�P>��2��P�
 Dt��)O9B�������L�#�X/e_ҋ�W焢��
Doa
�<����}�9[=� &6l����ţ�!���`��gjMҀ��v�0�^ylU��0Hv3/�Jg�MIt^%�)*�j^JF}�,D��(�kw�v��B�lAfo-�<Ђ���%k��SЪ2��Х�nNӴ���:O�1(��$m�
Fg�N���n����s�\kŊ�Oݞ�!�k1�q�Π;x!�E6E��=��OR,�`��b5��Q,H�}S�ˈb5�l�
�����1�Òm�M�"GR��)6&�Ԋ���n,jd�"�5���P�D`|���c�@j~"0��fc�.dQ��l2�t�8�>d�)�C�{�l�)� ݡ
endstream
endobj
32 0 obj
<<
/Filter /FlateDecode
/Length 638
>>
stream
H��Mk�0���>2�}CXh�ɡ��o��PHK����H�n$y���C-��X^�gf4��׈�v���fgF��j�\���a�1^�?����id4���dA�������k1�g���<Y����\��ŒAFǉ,c�v:׈��������D6[/���d֊�"�_�Q�wW�u�C�o��ˉ9 ��X����� �2���V�׈�Ό�z������A	�݊5�YFW�,��!��4�����l�?ȝ'�mSR��O:���g�e�-7�MKn$ìd���2��e|� {����
�����j�Y�H5��E�S�1gk���_�_^n}����o��nKN�^��Ém�.9]�����t�J�r���.�]Ӷ+�A�*��=e��uT)e M.�QPtz� Z�� 6ʩE�lF�h��*9j��2�+�E�y6��0^nזk���/��y�L��"���)V���=�4uᷔ{*D�z�_����0��"�ZУ0�V�W��*}��/Sgş�%��@��T���}�4m�6r0�z�V@
�>1�K�A�U^��뱔*��-�R�1P� �]�W�]y9�6��|��h�̳I%�z�W�t��Q��t�U���r)��7�Q[�<�0 ���
endstream
endobj
33 0 obj
<<
/Filter /FlateDecode
/Length 650
>>
stream
H��WMo�0��W�<�EQ� k�v��0�0�������H�M%��Y;m0�жb?>>�/�c�D����r���{��}��v��z�z����)0��w��@�x��!�=�?���{~]|�DAV};v��C��,_z�����}���	�c�q�8G�A����l����MD��C����ˍ�^��/�����W	]�y����c�}�'�������?����@h���s�K9�Ul"���	���H����f��5WӲ�&Ad��a��pB����PP�K�v��❣�2��\	�ٴ��ݓ^u9�BN�C�����5��n1ރ[�\����9��*d��w�5�f⥲�l��< `lH!��$���!h1Zr�LĜD�O"-e(�Ta�4�i�4�U,2�� ��]�9g���U�眩�23l�b���l43jKN��"Ʒw�U2����Jn�O���2�&��Fj�H��%��9k�n��+J����tIw��2澦2*������I*^�c�TQzV�7�Q��X�Q���Q�sԊ�����_w��d]o>g�׮���5\f�wZ��n��RX�^,^;d���_\Ba�<7r���ʟ8AWn�.��.V�i{�U;=�QWՀZ�l��I	S�9�m]J�[� >�!
endstream
endobj
34 0 obj
<<
/Filter /FlateDecode
/Length 718
>>
stream
H��WM��0��W�\ةf4�e(�$�z+�V�
�R����:#�IN�Dr�q<���͇ޜ:���5��{������$��ޚ|�iDp��'�����lɯa�3�֏��,��ؽ��W� �����AV.�w�A�_�/�1��C c��|�<?u���t��zΟa{�Z�!���[�������z�,��	䔉P�Ҡܖ0ɪO�d�f|��6�;:�g�C١u�������&h��h}�Z#�n�?+ �- ���U�,⨏���Z�Ӥv�d�C1��A4���XxCR������>_�1��J��M鞃�A�(��j���K#��rn��g9u_20p�!+D�l9����h��!�z�GF��$"���q �l 2���s5�q���H�QD(�vIrS$�0��Z��sQ^���_'�����YO`�����&G���>C��Py~�p���k<�A_T�E�h3�כ��ue�g���PZY�d��A�ʙ�䫢�ڨ����F�#Պr���:��ʧX�Q��F,����6i���q�t�� }2�YaT��iC"�k[W�����Y,s�?���J+͋ ���]�c��5q��+�zh��T�y����n��t�z�z"Z@�SX�ݡ����,��5��c��LF�;��Z�`#V)���wiݘ��d`�����r!֟���  �0��
endstream
endobj
35 0 obj
<<
/Filter /FlateDecode
/Length 615
>>
stream
H���M��0���:Vh����&�=�V��Th������3���rX�4�1;Az�H3�;����u2:ze�zX����y�@�����J���Yۤ���?���R�w	�k��b�G/ӯ�]���Y	 ��Ay�fQ���1��?�+sQ��)s�](Җ�}m�%j�Y�u��TzwxH�P�b����x�1w�I����n֔�Kp�A�=g봷E��p�&������"�]hsfx�֢NI����䲎���Q_~?�ʂ�U�إ��-l9ehy�[f�]ʨ�H"C*1ߧ+sWr�<� AgR���+K[�{��!4cUQ ����L$��2�.�������� �����yR�Rͩ���%�N(.�Uf��D���OE�h74�O
5���y�H��H����62��}.��Ug��	�s���tb��	�>�ޔ"'E��W#�/]}bI���F#1�$���A~]���{�ѡ-�	��樉���L7��C}�O�vHW+%�{�R�/V�Q&i��i��Vj �z�J	p^�T#Q�Jm9[)y���G{�RR�u�ReCVJn����m-�8�.F���`6;���`��榇�"���(]`�+tqTo �ۥ
endstream
endobj
36 0 obj
<<
/Filter /FlateDecode
/Length 669
>>
stream
H���M��0���9�X��e`g?�-̭�ThK����P����#-�q	a<����"�~�ΗI+og-�Ѓ�8[�Ut��:}�Z?�.?�����~��:�|������O��!��l�V4�O���uB�,���:�4�7�6�1}�^�ؐ�UȔ}fi�OwAi�|y�3��\>��<v��oHIl���"��4(�e���$m��fxE�5H������C��
F�:��!���%�W3!�}��p	�|nJ��4�����?�$���"�ievg>'��uJ�LO⃱
G��{������#h�
aA�W"��.�6ț8PY�+F�k�m�Β�i�h�6$��Ux1��\��	��������$@�T���f@\��F�
��4 ��H[F�֖V�e+�b\����Q������ÛVjA��.�J��}�g�3����γ��.��X����@�Q{�S])����-{׆�@B�e�2ʥ/�>s˙7��#a����\{��x�����֐�㥞�=�!wʍ���W�\�������U݄��F�?D���Q^4���By��ۅ��m{��WJn��R���r�T��D_��z)z�wX��Ms�^}z)��^�zNcFӸ��j�]>y�s̥ɑNX+, �+�yI]�#��L���ߵ� k��
endstream
endobj
3 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 4 0 R
/C2_0 13 0 R
/C2_1 21 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents [29 0 R 30 0 R 31 0 R 32 0 R 33 0 R 34 0 R 35 0 R 36 0 R]
/Parent 2 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [3 0 R]
/Count 1
>>
endobj
42 0 obj
<<
/Count 2
/First 37 0 R
/Last 37 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/Outlines 42 0 R
>>
endobj
41 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227171703Z)
>>
endobj
8 0 obj
<<
/Type /ObjStm
/N 21
/First 157
/Filter /FlateDecode
/Length 2658
>>
stream
x��Z�nG}�W���@`�/@`@�(�d�Ȼ 聱�Y$X���S5CGZr�,6�uq�/��u�ncM3��lB(&��c1EJơ��ס5�)��*J���θ`J+�xo*��2z�#�d��(��2�LM#V�,>F�`�7��lՀ��b�}��l���˛��G�����j��|y:��������|1O�?�[��������'�0v��4=�}�߭�����˳��8������������7&'7��\jգ��l~r��xk2����������oV�B5���|����?��V�+����i�au��9�o~Z|Z����ׯN���Q�s�|���:g������f������R_�SN�o����������%&:?�,?��TPo�\�wV�dnVכ5����e��������Bi}�EߧW�^��sx��#��@}�����6����k6gέ9O� U� U��
J�z9jQ0!fA�Ѥ���
|�ַ�X�H�K?,C�ڦ`rsxWM�T�dRF=�oTwjgt&�w.�$�jE}�; ;�,��Pejtv}�-!'���\x֒Z��X���1��Y&��L>�֣��s�;~+�-ql(qB�Y�r1��o�|���7V�Ÿ�uR�,!�^>�uzy���r�%�� +"Q>�|�^c}���6���>p,��̳�ڝ�t�K�h4�2���߀�*]�Å���`�B�N����H��£}O�0�6�;]�-ǫV��EI�";U���ze�
#�2�(K�0T����AI�9�U��$T�!DA:%I��)�@����ް���}Qs��(S�eK�@Ȱ�(<� �'.�hS��Z�3`u��M��j9��僳r�r���c���2�����b2�T�b��E"���D�Qi��!P�b����"�։(��oA�!"�Je��� `�V�� ^�T��.�YRk�����LEE�IߔUF��'uX���B`���T�sɲ�:({�^ $�>�)P�1�� ,�,�x����b�	�7ǂ��5�����hᶉ�&�!p��J,�B���!�XP�ղ��tXb'`/%-H�ݻ����$��D7�n��t-2,V\��_��|$�,{
��X�o��X �y��K�h
Y�L/�aq�c:��n���!��Ne9Z)\A���^P�0�aĸ]�WkT0`���؈����>�c���;�"�(4-��Jkf��vI�eqU�X���ʗxZ�P������d�S���1y�w9��p���`�<AJ�{���aK3b�PG���˟a��@�6D�)�"��c�EA��eT[w�]�D;�ЃY�-�f`}��ʆ��. ��76����I�� �w���L�z��!�QL;�ro�a��Zr��ދ�;�˹��c��Zr_�!;��}̝D�Ҍ�CH�ABZf��K7Y� ���q;���u۝H�E��xX�x��Ăi�ޥ��l;�%��'�5"��>�l��[6�s�ؖu�~�Nt��Af_þv��֎���!�k�yhX��z �y��{����H��p[�O�w��W�Na)c��s�0V�
��)Ж�d���HHD&�}��I�i��	y��\�y�$������x�+�8��m�iH�F�4�d��D���q5�,�piPS��*�~b�MAx����1����n���>������q��oW5�q
���|���3n7�����|=��)��e!�b��"r�<@�;xl)L|K:[���QҦ�x�7m�5Ҿ�g�{��swd�t?Q�>��9��1SRp,�)�����%GPLT8Ǩ���c��"�AP�1��D��.sk�c������e��d	��L�v�r"��C��dZ��.��IL��"�Uq��9�?�%��J��D�d�X8����֥��	 �d�D�1/'�������������㰋=P�'ѝ�;�C��["�0J>
�c��G<!N�L��3���@SNJ��}�Y�8�l��<��>���ki�a�e�0��ꀾ1{p���@M�>�'Oن{�5�����]��w����&��{���":�{	�����	&��_A��z�*��^���`p�C�|q�ۯ�̛���-ػ���{o��V���jÚ�&�E׫�������7�G��_�����W+T\���܄���uf�y~�@y�S[�׋��9ry��&I�#��R��J>B5>�x�e�r|��G��G��G��G(/+�k;�*�R<b�1�)���W���g���G9���C7���(��*q��T�#s-�����F�A���Uy�2GP�nQ)�G(y���R���6Y)n8�╀P�$��*����G(�LJ�F\��G��G(^*U����>��>�ƺ�]�~w��k��t���ޝ[wUy�7�.�׽�������ӗ?.��,��e��^�ם����0�}�.�ݧ�]t}t�>����rl�G9�2�T�]e��U��{�g�.����.a��4��&�5�I��W)P���<��P�|��O�*�'T��?C�|�*uO���83��oא�9I��j��+_<��1ݷ���`�O�?��կo�?��^�Pȡ�A�"��/֟� 6z����P�����G�k�}��Wa�G
endstream
endobj
43 0 obj
<<
/Size 44
/Root 1 0 R
/Info 41 0 R
/ID [<820C1A958D8B7D94161CBEDD213AA2DA> <00F4455B1AE8FAA902EE7842D7026339>]
/Type /XRef
/W [1 2 2]
/Filter /FlateDecode
/Index [0 44]
/Length 149
>>
stream
x�%�;
A����vt��y�LW1�@�(������@� �`�b��E74���0�&����**�	X(baψ%I�8k������o,Ѵ�cO�EGtm�E*�m�n'd�aE�3r��\2r}ĵ�苁�,L�Ǜ<���K
endstream
endobj
startxref
51818
%%EOF
