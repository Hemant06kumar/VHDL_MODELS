%PDF-1.7
%����
10 0 obj
<<
/Filter /FlateDecode
/Length 22
>>
stream
H�:�` ��4�Ai!@� �
endstream
endobj
11 0 obj
<<
/Filter /FlateDecode
/Length 2329
/Subtype /CIDFontType0C
>>
stream
H�|TkTSW�1$��2�c5Wｶ��/|��8���W($B��BA0�!A�^�E]�)Z+U�v��Ǭ�Z��9���27�Ϭ5k�����}���9{�Â�fA,ka�_D�E�e
�V�+C��i�b�˹�B�EE���E-p�0w}�v.�Z���y��5o���&�O�>��0��A�,w��2V�'�*�2�v��U����//�.\3�kgp�n���+�����3�v�3ZD�V���U��"�T��J�Z*YE�LN&f�U�R��*���\����L� Ub�/c�R	�V�%R�X�D�.����'!S����X��1��B��Q!g�đi
�R&U�Z�&ҦH�̈́Dz��,��C(�
��A!/���B�P$�¡/��fx@�we���c�����}V�Cv�[�[�4g������&���2��2����ٔi�T����`��<�	ho�B{��:�p1���F��b�������iP��Glj��س�`�AH�`QZpz�Q����Rc��)�ws=��Wt��e�;gS����G� .�,�<un����ֿ��JM�c�[4�n{�[�X_���w�_�����5�\�_�w��-�|	��a��\j� I�N�5�::��Nw���b�VAGS�UsR�J��Ф��yԵ"����7��П�U4��!�����x��Tfz�~_`zS~�⠽a���D�S&���>�)�ϡ�gђ��b�	yb�>$!A��+W��+�+}���W��9ǹ@�l��q����rK�+�����.$a�&��z��ꛤL���S+�aڃ�J�E`)��� �, � �^	�޸&^ >�h7:�}��f�K��� M��p8�k�:��\�� �~	/���޷	���)m*�{���_<�щ�u\��X8��gǚ��V�.&��,��B~��Sxc��ˀ���o5�'�`]<X�#kp���Ȯ�3����i?�#��'�*Q�z�@ 
����2�l�)mE�݉���q9�Q&��Gyԧ�שq�OP�aOr�e���X�3K����j��0�M��K�����O-��2�AW��x�%��.��َ#1Y�ͬ��w�����&�{���ϗ�`e=��FJ��G���6z:f��>fj�[��:�����'�Ƿ�t^�oe
�?\[1�j-	��e+cR#���1�қ�C���֑r�[@�wrO�{�τ]�9�i=�(b�*����&50��u�{-Ɗ���=�ƾ]ֿ�9�61/'����V7��X�`�}6��[�m����:4C[Տ�/��임V̖&���P���� �Y���B�]c;u�����[N�D*+�,u��ӱ�p-���I	� ����H�K�w�ζ���2�Y'����9U��o�tmBFj!��<��P�m��+��O �g�[@��e����ԜwY��h�{���*jJ[i��N�`���𔃱Xl��_!���30���m�[��
��>Q�gZ� DT��T��{�!]qD���c������z�ؖn)�x���>��+�y������b)��7�7D ��ՊD���$���9՟��_:�IJ��,�.ɰf�<Ҭ��#��Ui%I�����&-���Q��~���W] �}(1�0���֝������6S:�t@]���|���?%��uvk�+7]��۶M"�)�ä7<�����>&_o�)�o��(e����;Cz���9����ض� ��+�S�5o�xL��4�P�S����Җ�@����)M*;s#0��)���<�-!x�h����ET�HvI~��������T�d�$4\��Q���T�|;b6�2���˯�oS��$��Wf�ej2��p�&Jw ��įe�MB:�3��a�@n���&��`{[w�9t�)���¾y��3);u�Ԓv��m��c���`j��6"�#)�XtuP�n�%���eu�*F(�����o~��R��x��,,�v!�
�p�����v��ѵq����/����x
�x��z:�W�9vN^�:[�*�~�A�?���� �  �����}�JIB]pn�����<�cʔ�����Y�gv������w���X�����o�e�������V�W�W�tӁ��R�}jie|g^`����ϋ����[�[�\�tĀ��T�X� �bΦ����N������D��.������ 
�&�	�|��I����%���������F�_	��
��t�� nd�
endstream
endobj
12 0 obj
<<
/Filter /FlateDecode
/Length 308
>>
stream
H�\��j�0ໟb��!�k��1�Y��.��8�8Բ���߾�LH�>4�$�,ͱ1ڃxw�l�C��r8�7'.x�&JRPZ���-��F"��y�84����&'�fxګ�H�9�N�+<}���f�h<�Pנ��t���֍
��������-BJN�0rT8�N����*���F�Q�擒c�^~w�ʓP�i\/JRR��2V�zf�I鉔IY�:�8Wp.۰
֎�%�߆�˹rÕ��U�����:���Tf����xͲ�vܿ{iL�?xt]ޜ�K�N/=���-���D� Yɛ5
endstream
endobj
17 0 obj
<<
/Filter /FlateDecode
/Length 23743
/Length1 51240
/Type /Stream
>>
stream
x��	xTE�7^˽��t��%�$�EB,��!�$BB�fV�]P� 2�0����`DdQP\PP��'*���`r��U��,����|����CU�nݪSg�S��iB	!��LM�[���+���������E�TW�|������p��.B]�}g���"��@ 8��	�W ������ey��*�k4P�ȟU�\g�n�	a�E�3�&�{.��흑��L ��A��f��-�]��SBnS�:\\�W`r��1x޿�z�� �]��j���p���Ҋ����=c�ᾠ,oNe�N����ye�����B���vheEu�{1���>geUa�������SG)+6��㲋���������y�x��ןV6Q��yn����Lezg���O+݁�����"z|{�x��=#v�Y`P'`]�C9G�=}�͸3��]R�0�G�p��7�����O�Aw11�(��������@��TF?�F�E�E��9R�����Տ�2���:��"�t=-��IYJ��MdZk�^E����2]Or%\%I4ƯSD�_Aΐ2����Eo-f�"qd=2
����RD�"��U0��HN���� �H�,'��YAg�X�:J���� ���>�ǳU�5����p`�#�A?�ҡ�'ZI4�~��3A�**h~Tx�� �S8����q���xz��@x`������	��b`Y�\V��uY<f�S7)E7�'�������v7B��0�p�}����A��Wo'���2������Z��UR�-%��1�fE�DK~�B{�r�z^�.\C�pl�ߐ��rV��՗t"�R��2z��ΒJ�8I/X�@Hs��f��L��t#��� W[ �`��z�,`�";���+ތ�y�Z"г!�f		l�d�P)C1ƌ��s��h�y�V��V�b)Q�*^i. ��F�c�9	b~k��"$���ČC�{��]	�N��Yp�=D��c�s��F���S��d?fχ�灃"ش�·�K������)ŀ�{9Y�US�ԛ Et&����n���%��T�l�G)���ē\�J�a����
v��$J�vƞ�/����,#_��ӵX�M|A7�񐙃6�7 W�E�@ڃu�CE�s��0���1J�ӝ4��꿥�hO����6]C���N��s�ñ�x���t<y��.�o��r���,������t����5rP�[C7���-w��er�Č�\�u1c�r�*�'B�U�;|}!l��I]��Ӗa��$�^v��_����+ݯ���ﾋ�lD��i�/���x���ZXQ-���S�����:���,|�H2Z5dz3���چ��d"��*g��37bT�^I"�aw��V����	�F��MD��p�v ��nh[H��u��i�G@�h��]���D�G`*����E`���|)���N�)�$	�e�
��	�;%�H:v�r�R��|r��� �*�:!����1�>� K�Ÿ�[�(�?��t@�IV`��r���b̝�K\�������d:�X�?��J�d�,Xo5��xF7Hj�C_n�c��>O/�|�n�Ы$M- 0
ze�)9F��&�@k��`�HOܭ�o�}�M�u<�ez��4�,r\��e�~�����G>�s!���ϒ4�`'�7�N��0)�?L^ �ǳm�;����f솥� �P��!��uFw'���wo�]�� y��OPB_ �(���1J�'
��|�>����ДUx$w�� �`&#���cH>�(��c�/`2v�F��!h�\�� �i��(VMiƪ�r̓r5���O����_O��R21�}$�TC��A�3��)�� ;��yl&Z��᤟V��4�D����CR�W�44����`���	����	�U�m�-�m8Ȼr�����|��Y��*<���d;�������^���尒�(��{: ������)�)�#���sPF�%��@�?ё�ހq��4��睄��(��3�N"n�E�Q�h�O×mǳ\����7�u$���y�0��c��1+Z��K\��:��I���9�� ��K"��oT�-<�֑�e��FT�鬐{��g��ݶ�d[�\n���uD#�e�,�M�,�K$#���"����Y�<.�ܴ�8�q����MDdպ��E<պ�QRo D�z�^���6�_t�������V5���MW��a�Ǻ�6� ;����z>�_���n�N�p9wg�N1Wߧ�k]�p������^�藁3E��N�)�s�����R�)�D�%�>��K��<�^����`w/�Ǌ�߲0������$�kP'd�����W��y�u��	d�,�# qTOB��#�j^Q߅�b��u2Ƿ7�0�ݴ��(�[��G>��p��p��Ƙ��=Y��;ɛȿ��0f݅S%���Lm�a^Z��+w�� =Fw��)�0��zc�@x�h\���<'����P^�6�E����?�VLp:�H}��>�� F��I�Df�{�w|<�cX֓D;5�z$&��	0��;܋�ӀC�w �+�<e�Ѹ���69��VRk��<��'����P���hI��ǍX�hQDDyP�Di����d1�O}]�k%�Ed�	K�]�!�)8����b��9�a�%�\Hx��d��Ц=��y��f�������@�w?�% o{
`�� �7��$��ˈr�?�DLs���ܟ��ϔ�ԣ^{EM|E��<ة��EF�\H��(�"�(F�،��+�9��*޶Ш�7���6wY�$��A�j�^E���hQ{V���5�ho�}��yFy���x��He�h��¾G����3
���F�r,��Fl?�������ύ17�����x�p7�9�Ρs��޼�s`!��I	��b�ފ%^O�u`%��u7(���I�v�  ��H�ƾ��/�	��)VMĉ��e�h�|��3~�>v��x�i�"aӑ�����(=� ��E|fF�/��tB�6��+� ?�tQl�X�����f.��EL����#:��H�V��/�G A�]��=�#���ꈬv(p�	Z��D��د��-�a�LP��|���]�C2C\{�XZ��q&q@��<���8X�d�]�%�A���],芅�
b=�؈\����Țڑ���a��Y(����J�����/v�P2�����v�l��� p��A8�G��ב��	{5��F&6%
e(J,x��1]�<�:��`�����ĉ�P\{�74u�W
iœ��#}q�G�mx�k��^"�.x��+���#�O&o^#��3�Pd�٤F�^��٨�˜h������tj�G��^���??$f�B㷡���*)�E�0 |���;}�>$"#�V�m�:�b�ҫeB��#���5�nb�k����?Sf
��9�����[�y�z}82٘_��ú@SN� >�˙��h��̓���s�%Nk���ͫ��{f��d�w�(��^"��������x�P�}r�'��#�W�ޡģ�Gy<��� ���A��;>?��֏�w?������ /��.�{�"�ծ�j}E���:�lh}m�K��ky5�+�#���>@Fz���*��G���ǽ��"��O����?�H���������蓒�}~�"��)̕���x;�(�%�c�:8�C�PkX���m�Ǡ��!�M��C��c����8E|�#cp�+?	���Ke?��+���_8�RPGb���3�Į�;�L�K�m���?1��Ũn�����=��H)��(�v�?�U8n��g�����&��}_<���Q��"��&3�_�w,���"�!���p&�%��(1Rk܊����M U��2e��M��$�<$���TzpU��5p�wɂ����Ň�>�A��$w�~&*?Z?�_�ǘ�=20~�8�l�X�v)�v�]A8+�q����O�gX8$!�t��w��Ë�摊��8m<x����i��a�I��ė#q��#%Jd�~v�!S##��;IJ�����|>����5i��c�8��YtZ�~����#z��p봛��I�~߹�z�;3W�Nܯv�ϣ����O�᧽b�d�:�ipJ�mʴdtf�)�Ѝ��d�L��_�ƿ�i����Ε��Q�W��z�-�A6ܭ&v�A8�9�ED��DG����(9uȶ]��dj?��=���jb4�E���fƩL�S��g����85ɶ&Ǩ���~.{�졮�:�u޴�7��'�_O��|�����pm����8�\�~�zm5��H��jW����{�r�+��wq�?��������οM���7��ؠ�z�9�[��H�������r�R�����7�ё�U�������������^矄���:�H�~�~������_�R���������w�w���0�����oYշu�������:c�C}��=M�g7�WWE������Y�O��e����S[|Փ:?���:Q�ǀ�X ?j�G^x^=��߭��<a�r��h�����Ky>���sy��D�Y����u�g�zF�*�
���� �����&��������?��O}*����O�r�Ov���v�R�k�ً�N�;t�[�o��n/�۞���B�v�+ߪ�Ǳ��:���7o�U7�|S,���u��ǞW7��1��c���)�E���\�z�?��Gp���|]4_a�M��ۇ����*mU4_��+t�\��t��R���Η:��:_��I��|�����_�.�����0~�����y:���Y:�����������J���S�x�K����:��yEy�Z����uW˳yYw^��{�L��$���|��H�:/�y��05_�Ӊ]���t>M�Su>�.u����O>�'�fR �ˇâs������C�;x�γu���;�L���:K{�cu��<ӝ�NQG�i#Դ>*%D��Y�Sq��<O	���H�G$9�|D=s�,JR�����I���.��&���zzw��6���]�t��,�p^O]�e�·�������ޝ�� xPػ�:p������:�7���������G�	����xܻ����Њ᱖�j��WL;�W �U�Ĳ1v�ӎ�r7*=o�V{��6��-��`��:��n:��ϣ�'��)��?��y�����g/5bw���cxV�yg�w�l;�#��1�w�y��Ct���}P/�}
��A�x���øv�< �t� �$n�
v���������ߐ���U��q?Cv������Bv�(6�	�����
N�:���f;7�\jM�j �`�_���Ke�9�'vN�i��5���;?����?�	�G�/���ED�,c�yA�6����q��U��B{iD��|G��e�K�E��D�w-21s-������Q>@�ot�\�6���mE�*\|~�|~��"�(#;�>`��5+�B�+����o�!�_XOv�
�eK@�G��)W�&v��3�qN�ǯ\�^@����aCY��=��8��%�|���\'��XO`}2�lU/���<p��^�B:k�Z�)
\��io�Aަ�S�>���?�K�(e6�L�2§!�C�����(�V+�s�i���le�C.�t�#�#��e�	y�e�jx.���$�F���k�:����(%�Ǔ��x���L�u��+�|u�d����o~)ڇ!scEt��iV�d��E���YJ��Ĵ�T���E,_�oT�՝��M$����Ҁ��Ԭ.A�w�|Cob?�p�!��#��(VHc5���W}����華"�d4��ᐭ��.��P�r3Q��(f��P`�:�!!�:�$�����S/4AO���|;"q<K�r��L�K�������&�{��x���"��m%�����H����arcC<�XP`@pTW֯o� ^�tɒ���6l��.��W}����\�'�w2�v��5	�&�c&!J��66$����> (��������d�s;�k�����C��/}~��$r�]l���� ����6�G3�����J�6�mVn��2	�W|,��Z��<�!J� G@�X���9):pO}�)�Q���TGG��S�B�������h��eͬ�����'���/�s_�~�x��t���U)�����;��-���Gvh\���&���l�jG�5�ڒO���Ӆ�
�E^Ɩ@o��d;S(��NJˉ�A��Y�~`Kvb�e�_�}�9Hv0,a�8N�wD�ˍ����Y�R��J:��L1�Z]�Y��lu!�6w	
�E����a�]@����t���Ļމ#�F�S��8-�g���Y�|���t8·+����p�p�p�p�p�qd��Y��L%S�T6�:�g�F��m|��Mݦm3m3o�l�n�y�<M�fO󧕧է��MO���<m}��(9J�����rT=�55���I�%b<K��Tu�6�4�<�"�%D]�wӾ��$�
Ԣ"���d{@�� ��u�u�졟��?0sܠ�c��Y�j�ëV=������ի���f��������MO��4~�>G_�?�ϡ���t���i
�B�T�K+��
�u
�S��H����qh�<�(��pU88
�_t�н�������(�����_�#���(Q�o'r����jjHh�1Z��$��Iߺ��
�c�ne�i�]:��ֱc��A����G*i��_;��Kp���h�ݯ?0����5*R3�F�$(��ɏ�Z����yү u��I�+g�����X0�={N��a���-x8i���	�_�v�&Q��8Y{ z�����]]�u�e�o��ʹ�S]�Fms�S=ڷ#<04��=�G�Z�{�^|��!7n�S�o��`�Ѡ@Z��/���=i?�цhn^�U���3ޙQ���]lڲe��G�x�x�i�Su���c���k�3��n\���]�ʪ�w�~������wJ-b�zd�lI�p��}	�I����Tʗ[��J�̊�o��golN�!�|I�rV�@�g&FZh���$�yD?vQ�Aߍ����4-S;7�����g����[���ڝ�PW�b�ܡ��Xe8�ΗՑ徛M{�x	��HbJ>��ϗ<��O��vЫCH��6��z�]m:�sB̗Ԯ���S��=��矼c�w����_������ZB��;����4�~&�tuQ���:kx���{G��J]����ёa��o�I�DۅGw�x���6 �v��}�R����`�rb+����4R
lo�/x챗������Տ���h�A�h��Z�\}�Pt7�����{���~���G�<�&����Ν����}���Y}�L5���F3�x��*I*$�UNI�M���<��6x7�(#!K,���m��mfn�^}��S��%�I���Q$��pE��H]7�.�W] �o���Cl]n��o	����#�㡶�7!����A�M+D�b[z|�ɳ����w �Ɋ��l�����,~�7�}����t��%ݽm좹�-�?w;U�r���+6�D<����s>qz�+�>?���>�����[�ذ���)U�ԅ��l���������=l����:m���N�4<�f�*�|���*��稜�$�.�/��'�࢏3@h<�+�Y�~=Թ�S��SqB����*���O��6zUٴ�4��j���Ԣ��+�ezu����y�t�qUG�/�A�*;4�vV�Y��	^5O�� mlT����A�y��J,$��Ό�]�{�\!����fET���F0�9��'�{_��Ɖ�_��	��%k���l�^�+@U%*ߧ��D�tF� ��'D�Qen�>���E%����O<Kw�;�^r�4e.���Ѧl��vbV���Ʉ�T�}�&�O�m/K�C~F��"zR�}�&�uW��gHC3=��QA�Dó���)��)�ҡ�%{j���V�ɕH�̀�hU1�hѪ�X��ՌB���J��p+|����U-f�&_�Z�8�������@�^j���d�k�2cO0qJ�vu����
�>L�6�b����|7���ڇF�Ŋ/ ����̹��KϩQM
�w�']���x����u:�w%uVK]�rZg�c��'4�����/���Щ����G�yN,�7��wx6'�6�#Zm�������O����.Y�AM���%K�?�_�����3M�_��
V��\po��������ol��˰7{co��XW��?����l�u��|s�v	6�[�� Hkq�ؑ���yNbx�`���P�J�;&��'�p�yҎ����?u��ܧ����A7�JZN7����P ����7]C��X�eyd����Y��:��[L<���f� !�"�0����w��r������q�r�M���4Y?���������c~�i��o�!�zL�c�"��� ����^1ҧ:�V�Zz�p4��I��<٬��� �)>�)�=�TŎ6�g]Ꞧ�=q|������΃[�#6�D��j 6�h�6�2�h��
�U`��i��W]eBW��WDhҞw���F_aC�l���_���I�ޣ4��7���FYs��~J����/�'��v��7�=SO�:�҈��[�K�h�P`��o�M�߀����#�#�$�g��&�	�g��T��7�0`������!������L5�������O��Q�|xE-�$�$�I_�.��KpS2�}�Uv��@� �]J�c�\̳���3�j��J�0F��&Ɖ��g|�>�;T��)qV����f��|hy�3F$���[)���E5[-�4��C,]i����ҟ���-~�&��#�h��G G�xD�����������d�ُ�{�������k�J*su���L3iI��g̪FM̡�69H�ջ1z��Ae0�k01�`]MMX�i�e�L�k�4M�@g�bM��v�:TQ�(�?�p�|B��S��=��~��Z{���]�,u��.h����`�%��Dy��x�͑pp�k��+�mټl��-��������HZ/�4�A�BV�׿��4M��/Bn��.���EF��Gc�n�A�P_��3[���d�	WhП��s�?�'��荎��ì>�M�k�A~�M�"㻋X�����t,-n�Y�~F�#/��	qZM�p��t�{I'�7�/⨈�� ��W'?7e��f�uL�����=կo�S�H雇����G���>d���Q!����Oz�z7-y���Y�и#�O�w7����0�N.?����U�⭏L
��҄8�Z��������x�C�C~Cen�����B-u!��ty���7#�a��n�h�l,�I�����5�����;~�+�R���,�3"e0�75����}Ȑ�C'��k��}q���>�A���7���XN�h�Tq��L��I��5laU�&�Q���E�+\��nұj���_{�}��},8�!��wi)��/z�kS[�x�i:{��c�dl���*�#a\����F̂�K�y��Ư��,��������9����L�B����71pnʹ�����L#yO�2_�9��u�����o"CL�"V9�v^��H��_���Y5[�Sт�݆0
f�`��;y�j�UO��$��wu��w�G�Gn'��v�ݺ�gG����C��n��w��@���	w/��v�O���
��#C��y����瞻�O�~���@Z?�ؤ��sW������[YX����M�wL}q���;?4���nݲ����^s�@�ډĻ:��,|��eu�f�#%#Cl��!�3xKH0^fHo���7��T�v�5K�n�}���˗>�r�CK�7}�x�+_^~�`sl}=�{��.���}6'+�ӷ���S�׈װ�� =ѐ}(�su���=f'�B��_��-GD�`#Zj������"��ɱ镤=�7Yz�����[2�����C�)qPϞt �-�������Ƨ�r�:@�ݐ�J;��\m��w�>΃���� �QB.B�m�"2�;Ã����7~W}}��W/�J���ҥ�V-]���c#�ٰ&{�Q����������/|𾗞\�%����"���U�5Z��T[�K_]����Μu�[�k$�S��C�I�5Q]�h���3`��y%�3Sr??�/�XYɉI�O���y��G�/�kgS�Ҟ==pг� ڎڨK��Ԏ��o������#}!5;��jt5y�O;ne�L�5_�@��4"���R�H��䂰zg���"D6�t;�?�.���hϧ��n�cF���8~nmF�>Î�룔 Ϟ��j����V�koY�~�?ǎ�?���m�B�f�D�=�ў�ҥ��f�_qؠ�] k9/��V��ׇߵl��._�������ʞ�}�c�c6���꫓���٠7�}��7���Q��ة��ؘ���L��������w=b�Y!��R~1���i��q��8b"����h>��b/ʭ8�Az�A�S �X��J'�t|n潋W����]��������`�����i�شsZ��Bn�^2ֳ_d���v��89���
O����N�XM~Pr�!��LO2�"-�B�.-k,�e��4��^���v-Ob#.��c��U�"!�z�v�T����n�K4�5�&�c��.��k?alᤉ�^��?�������z�8��:�-���H�;W�� �b"�;j� �j'?��x��D��Z�c�F���R��W�����ș����>6pb�F�Br�|�2đ��ī�Z�)�o����o?<xx�����w�ix��a��"e��H[dZd^dYd]䳶���!kC�vX�qm���׆Eѻ��lJ[)�EkA�!�Y2zY��~����4:mГOF�O/�ߌJ9�_l��]=��M��+��L�6dxj��@7����Υ��Nп�e�ni:"�O%���/��d�M��� �d4,D:����՛�֯�Y��u�V�Y�n���}u��5~��w.|���w�ߪ���\�mڋ��-V�{D��`]���:5��#~��	~�3��H�[�Z����9��O�y�����s�=���W�6�+ˌ3lٚ�3�um��%�+Yg&��=ǘ�Y�L�~	hr�q��ɇ��;b9nB�B���'eV"Ο�;�;��I��xO���.�#�.G&ɤ��LG���8�Zt�,�}^�ރ����Y������;���2��#�~�t���n��咱w�'�F��9,DF�Ad=��
:�ڡ��>��~�������Ȕl~���ũ,ÚV!�'�1��Z�q�����6n{������bM�[�g�8�3���)�}���v)�����#{��(�[�z>*�H�~��f~��������ެ>���
�S��� q���V�����~mO���CNʏ+a��i�k���ЧL�}��7��#G}B?��i�}���z�M[K�y┎ʔ��f+=n�l46��kF.�ν�Bs���D�=��|��Oݻw7�-6��jl�O;v�|j� <�)ӈF
]= �6��`��	&D��qU�壪�FRL�\�B�ݘȎ�D�d�fEQY4c"��xT�Q�BS��U_ß��?m7~�U9Zl��J�A�n�XE��cYФ��&D��&A�C��-ɪ2n�9�c��X-f�7,}L$�C-ތ�-�F^o��Vy�j��N�igցwRB�N���>ᶮI3���z���1�A��:Hd�cbK1�YR}F�ƛs-|&ڊX	/RJԙ�B�Yl�:�|��ʧ��5���p ��[{���06Lbe�h��J�b�|���U*�����!���OG*��(u�����8qP���O�C��YR����i���t�r)d�C�r�R�5��s�$.H���
�Hk��J���
�Z�!�$�I��:g�K3k)6��Ɠ�w#��o���؂IJ4�B5S-1͢sM�g�f�V�Z�R�[���¢�c�>,T��W��z���Z�W��=h7eZӗM��E}8�B�{�c���ۋ�k ��J������,�`X�#8�؃��D\v_?_�`??�${;_�gYm:��;��a��Y}�9 �/��H����4(�y�����M�b�egf�9 ���կ��@G�#-`��U�+�LY��� �)b�ؑ���+'o(�c�H}�	�NG��ŵG�gdl�rR�h��K^e\^-$����P��j?�����֑T�(�Aɳ6J|��8�#3�p�hi��Z��
;IW��۴P��W������R�)Ȕ�%��!�62��!_4�"Е!� �FT7O�-�n�[(�������~&,[_�Gן9��;���}����k��f��H�+�n
�~փf���|�F� �	N��cB���Mi/ɒT5��P$�h�<�(�  ��?0h	�g�:ĬiEI�f���j����m��,���&�#���(~��-��&�E�J	�i��j�%����E�As{s�y��HK�e�^�� �ߩ���G|��h�'|޷�Ͳ����d��o�u L�{�?���:{�^G�-�`�-���܂[pn�-���܂[pn�-���܂�a���[p��	���ԯ�oAM%޿�D�wF��T4�է�~�U[%6R�ikď,�����X�i����	O�ײ���i�����*��zڔ8}�<mF�>#<mު_i�VI��O[#�|�=m3��Y�i���>���}�u�Y<m?R����s�Jf�8���p&���qN��L*����*�+�q����:KK�YbT�3����jVaA�5�pf��Zg~q^���jg^U����YY;��$�YPQ�WR���W^�[Q^�TQq��ªꒊrgBl��s�X<��.�(�B5X����rp\\�g��VW�V�UT�(�-/���]rOI\IyA����ʸ�������T9[P#8j��ٽ���9���bv�X�A{���24�9��������.[�+��DgMU^AaY^�=Ί��X���Ue%�R�]\XU��fT���8���<��aH/�YS��+�묄*0�bz.)��U�A�YS\�QD^~~EY%��5��^jH��=R�$��8�+�K�$�_[VX^�W#�)*)����r�3���f6d�CRRUXYUQP�_(������5���6b�����A�쒚��SV�YH��2D	���/؉q�J��~��cZ�#֌��rVB]R=�߰� h+��k<���.�(�����ڪr,X('T8�+b�յ�g�׈Cƥ0I�P~EyA��z�՚�Gy�+fJ+�4AyE�Pm�
�T�X���Y]���z�2`�ym��(�]T9�*�
oʶ�fneaQ�5�j��,o��_VQPRT"-������H�щ��W�jK��B��%3�%3J�VW�I�B��Z���S}�J���+m��$�y^ZZ0���ҹΒ6���
�7�ɱ�Q-�)t��"���B���U����)��>pF��)��x�h�nXk��Ĭ��f�
��`�8�*+������|�b��j��y��XX�V.X�����p�]�m�J���i���T�l�:��<g�� �/ށ�y���� c؋�����7�6K�i����"AԨg긌g��Ԝ	�Y)δlgfָ�i�)����l�G�8'��wg�#�3r&:ǥ:3&:Ǥe$�8Sr3�R���㲜ic3��RЗ�1"��䴌��$����LO���9��T���l�llJֈQ�MLJKO˙�LM��8S�4љ����6����,g�Y��S�#h3�2R��J��0D#�eN�J9*'�r����JLN��5&FP8,g9�XP	Δ�br����tgRZNvNVJ�X1VHgdƸ�BFwf$'植�p&���Ĥ��6�2"=1ml�39ql�Ȕ�E�0;-�F�d�d%��8�3SF��䘖�2"G���!�tI�q�)w܉��.��J�K��D�!)��g�]�'g\VN3)ҲSb��Yiق�Ԭq W�3�wB�Byz��D�ϭ��l��)��@�-���XXWʜ���a۞�m�G�J�#��p0��ظF�l����cx���%�����֍��p��
���+����dvI���8�*<�^u^)ì�Q�y��V�Lf��=+�J0evUI��3��U%�<Gq�稺��ʍ�WVW�*�UX:7c��y&)))GV�a]�/�f�ׇ�8gH�`�Z��JF ��$sI)!3H1�!Nҝ��&�x@��c��$aL��.$y��Ġ7��c|���R��d5㪖w��b�,�i%�h���#�16XfȑN�~'����Ę��[�qN̯��y�ٍx�%�a,F��$�T�{�\�_�Yg��C�����w��58��p/8�}��|/�����W�k���%1�Jr��Gf��{P�$'b�<��J��Kn%=�$���^�xu�s��g����BrX�������ʯ5��ʆ���jM��m�*�������'���/x.�H�)��I��I�ރ�
����Ep�)�Il-k�.��
=|͐��K{,�x�������#骐�����]a� ��ƣ�i/�I{q�H*��<��b�B*=ؽ�h���66-���J"����^p�/-��_�P����a����2��F>�ʧ�R�wo��e��5����[d"z*QW`�ZIg5��ik��F>����+�x�R>(��X�̖6P,=D�G2e��5G^�Um�Ҡ�V�0��vD�L�ӫ��[��1��GL3�q�K9%fc?�K<Rm��_��+9���f�����Z8�-�Q�o���E�Ö{8,l�b���1�*$1#�%>cLk;.�xI����������������
�Zt���H��@�.5��P�f�w�T�����<�y45��o{m͐����~E��Drzt_&�����Ř���"���6����B&s��/���D�e�G��x���cP*dZ�J筭�{~�Uy�K����@R*�U�J3��&�S��y%�͓�cخw��S�/yj��
�XX����(�uJڮw�\nFc�G�r^ɯx�*�*�������n�Lﾹ�)����6�-�*��#or.F6�}�1�{�F��6c��p�L�����������,<-���DLV�9k��J�q��I�Z�<����}�KO��j��Ң~�^�n����ZO�Z^���D����t�VK��=�[v�wG���9���h��RZ�=�gx4f���R�7��_x�_�j�g��x�ŢfI�")r�q$wb�q��!Of�g�k�����d<��WD$K�$�'�y�܍������D��K��D��Ny/��`|p��)�+�Ċ��8���M�5�3N�_*u'�E{$Ѩ�^f�Ƚ#�	ZJs�߲j[���^���.�Gy�&�/�M��&��Se;���T��RF��9��;�{'���-�(y6�͐<���K���ЄA�����9�
�R�gd��P�,�U��^��q-�v�X�,:���7��-�O8%�9�ɑ�I~/^�팔�6�ѝ��D)�qr�$�LHQ�3�ydV+����z�'˕�D�oʉ[[���:�+����HI���ِc
Ƨ5���&yᑭ�Ӱ{�&�[Iw��Qh���ⱩD)��\;D����DO=���Z�����f]��V�s�L�{1E�J���n�B�ܿc=����¼z��c��)k+_�>��w|��˻v[&K{J�P��,����])8��e�c�k���=�[G�-Qi��3����֑��Gʱe7�k�5��qf��<�c���\�,و�[�_o�a�n#7j��8݈������h�Lf˧-g������j���Y�gƍ���2OFb��H��N�3�Jy��̖�Od"������nȊ�nȪ�����+�WI}W#�*��d�o��g-20ޅ�ݠ�����P!��(/�h�x�&ִ� ����p���k1b&�;��o�C���%�-#�-g���¶��8�-�;�����v��ۃ����h�g���#{�C��/���~����iv�3�|B���e�+˕7�~Sy�s�[h��|���>�*�E��\�=M�m��Y�l���R!�w`	z�d?��hɩ�9�k^U�t�?����QUx�,ͫp�ɥy5�Hv)	����Ť���fg%I���zV�����Y�%��N�w���e=v\:����I��1٢�=͘T�Q(q�:F�}��)�����^ �1K��*9ԈIrin�/%�ٞ���� ���ķ݊�� ���\� ��6\���r�qo}b��x�]�=��\�|�NX�" �I9PV�tI�V��b9�bIYW"��c��sX�)R��'��˔���re��HY"-SX����u�2���.jRO��>Lf@���Q��R����'���������jl���_3Ľc2�6��Ʀ����2+�==��_��l��c�1������b��F��Zצc�rԯ W}�~B���;�#ՙ¬��ڳN,�ug��/�\,���,�˦�?��*�,v{ ��a��s;������a'�+�M���}ƾd߰��:'\�6�Cx��o��?�(��s�]|/⥼������J��o�[�������C����o�������_��x����O	T:(N���$(�aJ�2Z�T�+���J�R��(�����ʣ�&�	e��GٯT+Ǖ����y�}���A�N�Q�UE��v���I�T���j_u��RS�t5K�U���L�R��ާ>�.WV7�[���.u�z@�W��'�W�7�w����/�oԫ�u�h�f��-L�ݦ�k��!Z�6J��r���iZ�V�Uis������:m��Uۡ���i�h��c�K�Y�-�=�c���vE��5���l�3�:�����S�i�i�)�4ڔio�]�J�4]�=�g������]Xa��3V���ִ�鬰��7Qiz��}��W��M�ȺAbHG�]V�]��S�ץ9�Jԥ�9x�Nb[.�M�=C�ɨ���b-wځ�}�4�����b���)s�ψZ�ۊNַ�K��U�����7�T�͕�(9&Vx�h�\�A���-v{��������A9+iڍ:U���o�����sd��Ε=�e�${����9]֓܏��˽U�EO��'ȞY#��z��[Ԡr��.�W��񢦟��^.k���k$%�EM���S��:G�������̕��?��I��K)�e����^�y͆K�^�uLK� [��M��5��m��Ӆ�&��q�!1YÉ �y�YY��I{�ڗֵ�h�Ũ;�:Y_-)u��$+�����Va�Ji���?Jb%{r�5�IӺ��,��M/m�O%�����'��d�a�7���&�wV7�����tX�AH8W�K�aE*�D'���!��F=Gk���%g���Y�ת�����]���PΚ��ns��{=��^sC���m�ߨ{I����	w-�3݋�\=T�Mϡ(0�l�{z�w�!�����R�e���<�m�l<@�ܫ��0�$��M����Sb�J��n�~,K�G]����HfozK<m��Zi:�:VD�O�/Bl��J��C�9қ>'Y�!�*{�J?�"<-,g�ǃ	��2A�� k��@�'I$��p��i�&���v��v2ۖdA��Rm{�<�^D�}#}���}{�� �}{�Ɛ�����˼����VMhz���=�L�7�<n���h�2z���0����3Y�l�=-�����=�,QT�"n�ܕ�+�V|���6]�m��Q��O�Ft?�����XA�`�τ(��(h���D�ҷ�{�cz�~E��k��1ff~,�u`N֕Ű6�c�l4�d��d6��rV��E�!��=�6�'���Avr�fǑ���γ��'����c?2�+���=��#yw������Sy:��|
/�3y%�������a��o���.�����?�_�o�w���3�%��_���h�M	PB�0��r���W�(I�(%C�Q�R�)EJ�R�́=��T�)���e��OyF9�S^R�*o)�)+����+�5�Qe�Y�S��S�ƨ	�@u����V3���du�Z���5�<u����Z}Tݤ>��T���Ճ�a��zZ}]=���~�~�6�ߩ?���hVͮ��:i�Zw-V��\Z���ei���@��Uj���������m��]ۥ��h�����������������vU�n"&�$N�M���f���T�حg�z�oM�n�Qx`e;���y�]D�^U��W)�(����S��*"E̢�`c���?T���80Ӿ
Ɠ/5�I�v^xr��8ԫ�;)9�UA�V�G�_Q#�u�II���"<����p��*C�Sd�찂肆�8��>Q���N��~K���Re=�U�T�.Y紪'�z���d=M�~Y��'��Pߥ����i����ɑu���������nQ�u��e�rUHUs�A�;�.�ʥ����-�:=$뽒�\�> �]�~�g���DѪ�%Y��ɖ~V���2t�Q�J��7�z�Tũ���P���W	������[�e�����m��+��~�k%����lf���I�Z�maQt�"ΑN\XH�*θd�HX�&�gjC16`g�m㧥�m�V*�z�xEh$F9)�b-�rEbg�S-��4ii�����i���i��臊�����'�xe���Ai�"
}O�S`�!�8�l�^I���,$�~؛�F��"�� �T�K;���\����h����Vi�gT���}gS��x���� =�7�8��.p�7��t;��WjD�"�F�iʝ��l_���/�W�T�i�~�>�
�w���.���Z��WD��4�/�a?���"��^Up]�v�Dr�����o�����E��������-z�Z�Ԭ��i�.v�V ���﫹��.��@Y�p�A���]Ƴ�DD�W���K���~Zz�o����pa���i��.&<��q��J&��<M`�8X��z�W�h�VD�)"R���0���LF$Õ�*�%QȨ�$]d<�]�32�)��L�m�-��ْ�܋H&�|�����2��(�O�O���.f�1�m�F}Xc]�m,��gCX�2X��McE��U�9�~� [�ֱ�l+��v�}�񞑽�β��{�cv�}Ů�k���?���y��]yO��0��G�L>�O��y1/�5|_����|���{�~~����i�:?����/x����uEQ��]i�tR"��J��W���T%]�Rr�)J�2S�TfA�(˕���e��K٫P�#�I��M��C�3�K��r]%���� 5DS�����ju����R3��.u�Z���U��~�Au��NݨnUw���}�3�!����zV}K}O�X��~�^Q����̚��uМZW-FK�jôdm�����&kӵb�\���i�����ڣ�&�	m��G�������*��>���;���B*��K0��1Ƙ�(�*T�UE 0�X`AeE�)&�P�b�1!
Q0Q��	�Q0U9T�P�S�C)�rQ)U	�	Ƅ�޹�@+O�L������ivvfv�3��s�Hs�%�99i���\��G:"��[�.f1f0�e�L6��dcX�Ȧ�\��
X1+e��RV	��Ul-[�6�Z���`{�>v�bG�qv��a��%v�]c7�m���˖�&����(9[/O���3e��&!i�j�/ ���.rbJ�Z�g`���y�nޣ�z;!�_��@ʩ ����:��î��{	D̓�W�
I���{�mYw����wԻ���!2I?H���H:&P���-㽚({�%ث���ثA��xۚ�T�<����������v[WR��ޥ�~�~���޸T����oI�����6��=q�?� ���)ѳ�+�Q��Ǡ�{�w��X��N̏m����h&�s�̈́��s��JF��c����P��P�u����[��o��>h!~�����O�V�K���S��5��H:YE�IƐud�!�d'�N��Ur�����)YB��ϫ�8�wRAΓ��5� ��k:�'�r�|J�Mn�;�;�.���4JmRO=�Jާ�t0��f���O�P�E�!ͦ/��������5�+�Im�*;��TRv+�iHiTiXiR���M��2��TDYS���_�^w����C��Y�j�Ǿ|�`s�BVΖ�j���a5l#���X=k`�����Vv��dm����Y�d�X��c�!{r��)�G�c�y�<EΕ���X.��K�J�uy���y=`�\+o�w�{�}���|D>.������K���|C�%�H�G�hZtP4+:":*�����MH�PX X� TEWDWG��ݓ��f�V�v�.�^�~����(�K� �-zp 6���	�;��$ �pL8��ؐ���pc��
7+��ZV��Y��XQl��;6+,�X[	X�ll���F@3�%�;Ǔ�6�9�E@{�#�	�[�.B�0 � =Q��d�F`�Tr S �J�R�+���`vP�N�U��
hEلe�)� ; { �  0+G��F��rI��\Sn �M�s�8n�� ��g�|a����$�� 39葃y	-r�3��ȫ�
�����f��o�;����A��1菃��i~�_���U���;�SAw*�N�TGMW���t�/D���T�lB����LT��" hO]�����xt��TAsj��S��uj�ڠ��TЙ�h��TЛ
zSAo*�Mmt��9�^��@w��hO�i�;t���4Н��r���-W��
�b�T[�-�*�׵U�Zm��I�նi;�=�>�vH;��Nig���%�vM���։ѹn�i� =K��ҳ���$}�>S���%�}�^�W�+���:}��Yߪo�w�{���A��~T?��������U��~S�cH�lh�c�C��Ɠ�hc�1��l�0f�F�1�Xh�ˍjc��ƨ16[�:��h0�f��h5�'�6�q�h7:�N��e�͘i���af��̑�3ǜhN1s�<��,6K�E�R��|�\e�5כ��Zs����c�3���#�q�y�<o^2�����m�X�[��f����(+�oM��Y3��V�Ub-�[V���Zm��6X����vk����o�[G��i�u��l]��[7�;�d˶f;v�=�j?i�������{��o�s�v��ܮ�W�k�{��Ů�����n�[�V��}�n����v���o�]N؉9��9N�3��qr���'�'P (��:�x����:��������:�x����:�x�s ���:��y ��+�k �b��Ku��]�b�r��An�;��f���I�4w�;�-tK��b�­rW���u�w������r���݃�a��{�=�u/��ݫ�u��{Ǔ<��<�K�����F{�	�do�7�������B��[�U{+�5^������y�^���5{-^�w�;�y缋^���uz����pj,�H�R3R3S���~���+� oB����j���y���@^�k�����ھ�`;��>�ߧ�����x�azSBz%�W&�����[������zG#�؆޹_~"��^�Q~��H_W�A�j
�~<Q���r�K�w-�~h
�@?���]WR��ޟ��	�s_dv2��O��x��5�}V���!��x����Z����?>�ފyjy|���6:�с�DO��LS����&� �p׉Z��f����9����G�]��iP˽��
�d3K�<�����Pf��,�ttJVW��1O~B�@]!I�0n<d�N���2�&��z/'ў��������!�Mf�xm�w$������{�L�{|xے�X�9��`�� ���l�E��bBW#NqԢ�	y
���wZ�y*�|����	Xׄ����_��<�jӗ`9K0=�1}2晜�'�0�8�����ҞDx3�f|�v',�^�}���j*�ڀ.���3�
�<���'�I^��Z���0OUBz=��'�>�j0���<yF����{�,,'�m@ހ<�,�!� ��<�'ks2}�چ�<�W�< +R�+�ӓ�ջ�[ɡ�S��w���'���>������<��ȟG^��y�
��o��>PN�� oA��g��A>y�^�	�ȧ"�|`�����E�=(s0�4E�)E>��")�{�1�|�%�K����Cp��ʐ���;�y0n{��&�ː�!
�<���2�\Op�'	Z~9E2�3�}�K�2�Ԓ�K��9B��e�8�N��]���M�2y�~?��~��{|:�ސT:P�%���\i<͑&H��\i�4��������^����ZO+Co�6њл��t}JjJ*ݐ2 �	���7Sޤ�)R���l*��jX���bo�]l#�Dw��l3݃_~��V�^�}��6�ׂ}��`���EڬV��O�Q[�,�� �'�%�0:+㲞����pW�x�+�"�����W � 7 ��&$��p�H��"���Q X��I0��C3bGO����9�.�yX|ŧt���X{�6Ď��b/`�ػ88�߂(=�_�(��.@]�W�ɣ�N��[��O�`k�L¿�����P[�lEX���|Q쑢�����@D�&+�RC6�Ցz�@I3i?:FN�6r�\$����a��hͤ��H:��Љt
ͥy���R��.���u������&ZK��t����?�B�s��?��-�W~Z��=��,��Ǧ�I(a�%�XKJ`�$�L�]3 � �ɪ0���r8�=}Հ� �'vn$��b����å߂x;�x	�Yғ߷Ϟ�%��NG�q��1�s
�}�Ÿ�r���
DsvG~���,e����?����~�'%��F�2�(�=;{�{�+�@N}6$ƅb\h!ƅb\��-ĸ�Z�q��XV�G��>�ĕD�g��͛�l>�0o�+K����e/����Ye�e�I>$�!E���[w.��W旖��
�s9ր�����o��SP�{� ���8Ƃ��+$��?6��#ɴx���xI�C�⿋=����(Fz<v@yp�Ǐ���a\�뤸^%S�h)Q�ɀ�:s�[&�\���v ���wþG$������� �O��?��$�g��0�V&�i�X�('/;�����K��ɯ�kB"�d)˟���g�s�y>�������������K����_���_�o�7����Ͽ������������=�#�3�W�/��V~��/���r��rW�-���?Ƈ�?����R0�
X������X�Hd6y�O�_�_�_������K�2��+��������[�m�m�]�}���?��W~�|����?ʧ�/��׹����`�G�	ѯ�0���p1xdI���Z�D�����ڱ��� bi���sy�煼���异W�j����k�:��o�y-����>��Un+�J�rU��\�1���.���o˟��>�v̛�ħ#�I�IP�wq����4���p�9��3�������4��Lw)��QE#����%�Qa[ӱ�|B��[��gH�~c�CdyS��=�;����kn�����ʿ�k
endstream
endobj
20 0 obj
<<
/Filter /FlateDecode
/Length 478
>>
stream
H�\��n�@�_�\��-YH)�/�Du� �.Rh�/��]vV�Q�0qf>�Pԇ�a*>���B�a샿M��y:��0���ݒU���LE4��_�y�ݎ����m	zz駓�F�{�}�=���Q����_��PIUE�?��h���H��C���9z�&~=fO2i�cL���m�C;^<��xT�k�Q����[����iCW�z�e��/P�;����B�`((�<LbD�W(�OaDh(�%�,�����T��\q�t��H$"iűjͱjñj˱jǱj�H$�5���~� u�������K��vS�b��U��U��U��Ul���YË��m����nxi���l�$"Y�0�d��������a� �Cj��p<.cEj��"��ptn�V2�޺��7�s�{q�Ӈ&m�����?�E�4��t�` {�=
endstream
endobj
25 0 obj
<<
/Filter /FlateDecode
/Length 14674
/Length1 35052
/Type /Stream
>>
stream
x��}xTյ��g�s&�B!�W	B��~���$$�2�L�d�̄���FE�Ԧ-UJ�"ET���������Zk�U���"��Z.�3��^��d���~�~�e6{�}��{��^{��3�3�z ��5sf���g>gl�k���UP8�;�*���Op�UVZ���)c�KQ�bVł�Og�=�ح/��^Z1*�ތ��2����&w����i������Yt,zl8cC@�[k[ꚮ;ic�g���:w��9�X�{�7���6���p1�X^�u{bL���B��z b�?�ރ�!�M�5?{�g�1���獾���_���p�i�{MK���7����������gV#nK[|�`�&v�Vַ��-��4���� �Yҕr���b�5ݧ���a���#΄����N�]L%�Z��~�&s h�~��<���(ET�1ΰLb]
��r%�z֢���<�4ƴ1�p�j]�oY����X����~�2Bo��
��Ɏe���b�PHO2��vG�p9��ާ�_g���2��}��w�A,��o���Z��W��yv-��=�l=�e��-�v���y�UQ�7���z������C��}�	��l![͖��ȷ����M°� c���Qt�+v5kC�%h��U��f���/G�uK�`�|�AV����<��d1�����i�^>�T��UQi$�R>���3���O�=��l��#1H��N���H�pZ:)�.n�)��-7۩�d�|�RXi
$��Q��d9zt�:`Ȓj��
j���ЋL0���%�βX��f�ۏt�r�w,2���Vȶ#TGr$�sp;OכP��`n�y$�X��ȋ����y?8f���l$d�R��I�Ss���Y#Vg�٠��I�Q�H%.U�6��`I�qqS�Q|����,��m�,�V��V6�c�"@��/)���_�%mXZ�ѐ����}H�hK���g��"�4�it�r��6ǃ�\G+l}I�mUw�R�W`�|�ٛ���Q���vBf=LB~�� �~������V�hhx3Kd׳�d�SZ�� W����B�2��֠�\h?	+�iP�p#R=�c?�L�4�0Ul��;���*��e��4zj��k Y=�8ڊ4R��*���gs�X���S�D�S��|Rw���?� ���E��g����J,)3��~?����y�+�G��3͗� >����z�k���_�K|�6�s�#1b1��8���>������%H>�����B>�/��(�0���Q�U���$gԗ(�S����:��#��w�w1���Pw���f��c����i�0��У�y�!s��dh����Ǔ�=�6r'�s,py]yw'f���r?����������[��j�K/�n?Z�W�^+�|r5�3;��\�U���ZXK3��4�m*�I��r�p�W����� m�A\���bN��+}O�豍�{F��L+������oZvCi5R+v���a��l0I�e%HIh}=��U������J��g?�1�C���#�w�`���E7��'��@��&B�ڒ���#m�7�~Й����܇�fJ��#��X�7��7��6��vA��(��x^��y���ҽ�.~K'�'j�	ӕ~�A9��1���p5�Gʳ3��v=h+w�j���(� �&}P.�Q�A��<��lj33��Pz����D�y"�2���ꠥ<��߃u�a-̆v����`�:�;p݁��q���χ�i���S͆�l�V�$����?�>���bd�߆ ����O�'������������f�>�Ѿ��T�`���hv��F��ɧH�H�Q�mM�l��-AZ���a����J֨U4f�-���O�8o������f�s�^����V�n=R%�D�W�<hY�<�ǁ�r��緁v��X��cC�B�_�����R=���A��s����]vSM��~��`��V��d��Uc��P?we�Fx��A-f<�j3aG#�Yv���,^�4�O�e���}I��<��χA��H���	�iR6|n���F)r�&�y,\o�,@MoV�'�ʖ��:�����n(�y("�,�5�� ��y�Z �����۳�C�%K�s8�ꚣ#�CX�Q�����֬E�s�X
��<��b*�r�J/(3ESQ�뢩�ET�0G�h_��#}��2.���d�̀�O���N9Z���DFV�Y�-��lEtV�%u��}{��Zs\�2���=��p%�Ͽr������U��#n�}���m�7�g���0s�*����^������/���s�您�:�u�����h?�5�)�םo>���r�R�%4��\i�6_2��W�ͯx<Q.�]/�e�Y���	���K�Q6��J������s�>�i>����v��7�I=��p+3�|�@g�!�k�i���`���H��"��[�n�
|���&�T##e�(
[�`m�Qz�=��l�����X���]�Q�Y��n��2��n�x2�`_b��U�Ҡt�u���k�3qMÊ��q�!�_���a�J���SC�E�A9�� ���V?^�6�6���b��t�sΈ���c��3�F ��$�f$o���c�|�)�(�.?R�Yi�9vK��F�C)kz���g���ՠF��߉�����H�j�N<h8�!G�|�+������2�R��]I'R��Q�u#�U�k�Z��p��@{&N���|����s��������5iQ���H][���{v�q�rt�{y�,������LY)ܺ?������Bf��D���$̼�N���Z�YIf�dF�Y�S��j�v����G�S��_Nt�n�о�)I�.,�cN;0��>�����:ExƎ��8�Z���j���,���[7+e�=�l��d�eԆ�o�/���'�?�O�{,������GX�Κ��RR�KX�S��J���%Yo���}8���U)�G�_���&<���&%ņS��Kd�'�v�tR,:�Δw�5ħ~��{$\eL��~N�֋R��>!<�,�ԩ��U�_ßN��H:Κ���NFz	�t��v<�w|���6�2��5�ɽEz�шa7��&x�X�JC�r��n�2<j*0u��V�"�>������~���:ۏ5U�~�}bڌe�@u��D�.F�4>�g�-��܇�M[�60���:q��?"����6&��lP���@�2g�X���+��Ԩ�m'y&hCD7���pbꉽj��pȶ���Ȗ���X�A��+1�#��2�� �=n�ڼ�\�>	:��� �GCځ�__��h9��*�@s<(������+��X�l8IF��ʣ����� ��4���D`G(��+|>�W�&,�Kh)Ď��;��-I-o�3��H��W������y)Hy$v�
����uH��x)�i�U����߁��Z1����r2��
�E��g�<������lQ���S�_��C����w�H��
~�[r	�����m�h!�^Ng�<����vm`EUa/��l�K�B�/)q>�=�z�y���?����ʍ���V�6`����B|�k�-TJ�ӾB>~�+N��e�YT���k��#���N��%�,�����(�T~.O��ncL\� �$�3���y�{G���J���ˮ��3��W竽{��M5��������� |E��B��ދ\g�J�c_#zA�G�X������}>���y%<}�z,,OhU�1���1̘�:>�l��V���ȪF�w���^|��Gb}b��);mg��J;�����N���`����Cp�%Y �gh�>��F���r��ҳ�d�ׂ|�<�����c�/�9B��������k�5���^�Ap��׏�yJ���u��e�5v�QG�|�7���2Bo�s1i��RO>;�#�o%���z����؋N'��Sn?�c���}:zj��3�[�ɷ�3���Gj���Y�RNp��"���s���B�,˕p@I/�ȝ_�zi�Y]n]	�Vv��Z��P��J�->��? �c�郏]��Ys˪\�+,��./ ��
Ey4��T'=���_����z�]	w�|W�w�HvXِ<b�g�O?#�:'~~Nzr�v���,q0G<�&��yā6����ڣ+���b_O�)��������i7���M�S�yN}x�b��M����dh��ݹ�O2�.S�8G��%zp���):z=7�>��<��Y�Gyb�s�+�s������~N���z�溜��]Sl5�wL����	�����{��{��=��{�Ħqwm�vw���wn|F���X�m|Flܠ�q{�v�2qG�z{������m}ĭ��-m�fS�z7�7��6xč=�mb�G\_!���r�:4X�#֦�5@��զXe�`���&��fk~S\�-ZP۲^�RDs�3Z�)��iMψ�jcC�ָL4�+W��Y�h���z����:\�<�#զ
o���զp��Mq�G,�*I[j���Ē�xdmq��J�Xm�)����pj�	��)��'k�mb~Y�6?Y�%�RS���h%mb�G�b�)���洉��b�91뜘�^��
׋��bF�ȋW��b��xm�)�NqjS����<��6�ML���&��6��bb�:a|�6a��Ƨ�qcS�qs��1I��1&I�\���x���"E������.�RD6P٩bdV�6��yX�͍U�FtײE�a��n��xmDw1�0w��8mx�~�o�]�f�ú��sEƐ-c�H�%}��I��DZ�$--Gr��M.�]c��~I���"�TS@�9���׷���6bվ}��=E_��>1ݵ>����i���$z�� ��&zMIDO���<'z�Ą-�H@mB��_�u_/�q_%��L�Ta8�kF�pvq��8-����$t@B�!R�XU�b5=N�y�AU��a�r��j�J7M�
<U������#�W؈��� >����=�v]+��%l)�N�5C�� ǰ���㌰�n���V��gQ7�r5�LdY[������8��ml�xE�B5�+��W��[Nh
"����w��,�3<�y:b���#VSp}���I�Z����Z�b����uP��{�go���[�6��-�sv-W���I�����α�������� �͎��v�Eu9���㴲T�N�Ύ���^�����na��(j�������u��B��b�v���w{S{K�����ENd'�q����(Ǎ�i�0�q�PX�٦�k�:X�\C=��#<F�VT6��SW��c����3qPb���A�*;����lsğ�¯������+>�,N�{b���1	�^>�2h���r�h2��C��͵����q�B���@�`/�&��`����t55.���p���S��']�r�qE��<Nm�ԓ9G����Ł���(<;�#A��#A�����i�o��|Yny������J�2M�2���;�ʣ�G�~��E\|w�L1JL��f��R��7��fqG��-�G⾘�cw�G�Θ}���_�C1O��]Ɩ�=WY��PÆ��ԏJ�(���������?=hB�k���F����=_UR\iP_7v��*�^&���S_�j���#G�s�'�������;;�o�����z��ncmB}��߷g��&���Bk9rO�9u�T��/O�N��],1��I��齒��䌟����[m����.�<\�����۷o^p_��#�D��{�Ió�3�ڳ���2V^>��Bp��;���גD�������<(z�,Y�ILvf�)�ɹ��:uRr��c�Y61l�)�	=��$s�g���&z�!�{���}��o�d����k�����Q<�T�����j>����|�2���Çw"K���*u6��d�XQ}��CEl���w�������w���;23��d#�������G-��<i�,��$�J<Y��	�������7�x�����˖^{��e~��W��K.��w���F�[�܉G�����J~ۓ������OͿ��_�-;����e%<�sx��K�7˹V.�=�M,�uc�s{q1��]�P��'k,��pl�ѣ���=��_�j�� ���R��+��<��t�����7?����ײ�%g&�K���Yc6��8c�d�a���N�$G�J�D�I�S`�i��JIy������7���_������X2T�N|�nN֛����b�����O�M�-�����TN��a5�x�#MvpS�֬iX�fM���Ӽ�����̏�=O��'O�l����4�E�/H/�i�Ç3�F���2s��DlK��w[��&3g/HvJ�%�>v4�2JZ�x�KZg��\Ϋz���-�;#���{�>���Scň������������7�O��yG`̡�'�ӺJ�s`jL��K����9S����IkS�9֯Z�~g�Xj�s`?��/9~�#9)mܰ��G���d����2��䔼\��q� 7lg�rG���Q2c2c3�2��Ff�������F��J��9 35s`�kؠ!C{-�aW0PI归������6ƍ���?ZU�y�Y���><�=�����u+��3��O�]�O�;n�Ĳ����-?�����M�<u�ĩi=2vn�yp t�3�z����dW�h�6�D��25l:�	=ⓤAÞs,�;33d�\/����8�@�q~�ySт�_��<��o������s�?������������5�5%��`I��K#�띦'H�K�P���q��*�����f����2�����#��,SR�IYycf�-�u>)%}���2=���uM�����t�[�w��S�
J����R�J{�D῜.���r��.���r��.���r��.���r��.���r��.��3���t9]:ѳ�d��װ���,wVYa*k�˂���ը����:��6���Ⱦk��l �e���~��c���X&�/Wcqw$n�]���̴�
�qε˂��ը��R�vYg�0�����]v���'�r��F?���O���7��]�j2]9�G�qU�u�7A��ݔ�*j��v�56��e������Wy=�q���zws�7�r����fWKkucC���kr74��T���y�f�+���Y��|ͮ��1��^V���v�Z_3����`�e�Q�W�f|��o��_��n�G�nX�0����]��R�2������Τޒ')WDװ����6�Vgf����qq����eQ��-n�%?qq���]]Fn ������6��+]�ڮT��ʼ��� i��~/ƪ󻛃^O�����C{Y����n^�j�|���:���0J��-��^{"�55��4�����hi�5,�T��	b�;��4�14X���m����چF�x��H\���j�<-�8�{[�>Ok���x XCuk�K<tꐅY�il�HNV7�}�A0��`$��-U�lk �8Y�&/IM��ϊ#K�9��w���n ���]��́l�Tt�V����ta9���f襎�+��rZ�Wxk�c�&)��5{���qq��rW�VyIˊ���4����������aV�+P�P�^[k`F��$��v�w5��ދ��
�m�ֺ1P��T��&�ZI���i�m���n��P Q��C�[�����_��n?��ꚉ��Ƶ-��IZ��D�G��@ב,��X
s7F�B��楃"Xln\�j�d����%����ʔs^"^؝�`���	��"k1M��p�ɥ�Fj����	�`5I���)�*_C�1� V���҂%�n��
K~P�21�� Eosg�`���Z�"-��:��4K�K�l n+��NN���(=�K�a��f���a-�͇�Ƿ7�NC�i�Eoc�djv�kfiI���tf墼�BWQ����taQAa�+-��iY�EE��KT�Т<��r��t�+�d�knQIA���������UZ�*�WV\T\QɌ�E%�\��WRZ�*.�WT	�����&UTX!��+,�1�y�E�E���\3�*K$͙ ��*�+�,���8��U������4
@���df9F)�W!@hFi���Y�+�Щ�,Wey^AἼ�Y��R�\�&��4\�e��y�Ů��ʊ��¼y���ά��yRGJ
�*�JK\��%/������(�+���*ț�7���c���C�ì���,WEY�"Y���gTRK��(&vg��T�_ څ����.�! @�� �H��+�T��WFXYTTQ���+/��,�,/�r>�Cʸ ���Wb�+�H�.����m
�A�B�qA[XW�oKPڶ��-�H���Yd���	�j�µpT�=ce��cy���%��,��J���nd�_�*/�`@���t&��ұ6��}/�n�`�i�nD�@���*�!���e��!g�r��oXgo�~{��*��+�~o�;U�*o��l�����8ihF�d�N�	N�Р���{ 8b�lW��|��2?k`u����c5,�6iJ�h�b�hdd?���p��-b�h��R�񞋕Gh�΋�}Vz�2����V��A[7��QKʒ�T�[�53������6����J���H
�ЪY��C_ZH��#�9�c�ЉB����H����R�%]�ք�6^'ӟS{����>�|�������I�lz�[�W���ȣH*�wj[@��b��K�y�̨��z
�ׅ�#��'�r��G���V���d�K�.6��q7J�<_hoq���h���Oذ�dn���z7�jiu%p>��7�"%+#zMD��v-��T�媣Q��=D��j��Ѭ�l/�����Կ�^�>P�3�@Va�Rck:L3H\t^n��!i���)��lZ�VZ����̹i-�k���A�-�e�5��&����~j��m-;�c�)$�A����:��@Fi%>;��A�5�r� Ն�����T�Z�����d��!��f�-Q����UZܶ���fG��h>�sݱ~��5rdE�E^�E���`�n���y�/-uXs�-�v���V�>�����PK�ٖ�5���#�����R/$
F�D�q��%�3TCc{����ɴ:+�^�q>�s�:4p�'��L�^�Nm�k��> ���dv�3U��a[��ayr�%��G;�˞�&�z��-۬%~k�H�ٝ4u��R'k#�7��k���h�����,�ũ�^��1��V޿�(��ZA�M��y�S9_�Qڨ��]8)�C�d=���誟�7���<�,�Mst1.�I����b<f���H�.�����M��1��e��M�]�k�;o�XMRy��E�Ŵ��]{���]7-�ڬ�S�e���u���^�X�چ�hL�dA{���[��]�M���=�ϗ^1���]t�<zɢ��^,�.��em�EF�+��JZ�9�G�l���]�$�U^Q2�h�� ~�Gg�-d�+����E+���wx�����^#A{_��hJ��W�S�Jp'�)�]%[�x����y\�B�Rh��w!���<���i��,)�ҋ�]6�r@I{10������\�/-ٷ�U����ٲ�h���B���!_״ ��<��h���*i��~���J�;F��U��l��A�]��EDO�E����3mN�HG���9ӝ�.���*H�y$��m	�0��,�ā5G3p-�ز�,���B�Ti��"	�<�_�:��g��,�r�l[�.zmra����E�.���J��<����,�0/bGH�<�C)��OuR�R�ő��Q�2��%�Mr^@#�F*.*I�Z�ٹ�u�G�E�����u�X��E�e�E$�[�M��-�(����Q��|�Zh�T鮳�
��wHa�@�gD�c�K�ٝ��R������b!�ʣ���ha&��y6��,,<�l�,�p�Y��un�m|�E+<v�, {*�9��h��Z���Z�w�}M���;wt���FǟY���FG��Em�����Z��ڳ:�<�1��v��)ي�;��p�a�n�l�z(N�b�@$*��_$2YM�{�ul��� �kI�j��Jˊ/�-����v��'���QVS9hG&R�V��į�r*�w9U}��e�&��i�[�u�j �x2ۦ�g��Y�N�����z��Ij�Y�8T�.�s�=���jr�8�-^��n�7�_��Z
�aJ(d��+�1��c
�΄r��F�(mW��|��C�w��1�^�����Q��_S_C�u���T?@������'����q�q�1�0S����b$�Y�ɒcƱ��S��,�dn�����Y�od���ޕ����s����`3���4!��VI���xEy>��G�����,��b����K����b�*����؊����|���� �ݴ�i�l�1��;����(��ǒ3�%��l�v,�
wU�����}�����[����}�N������S�Y�)��?KLcI˕��m\���M�C���9�3X*�h����,���ԑz�z�B�Qݠ�B6$�"	��l��\���r=Z�r�(Ű�q<dZ;�o��G`{�bj�h�&t^
]��,s�Ю����Mn��&)����U��ӂQ��rH��,���7�7AGH�m]����W��Z���~�����芡�PR�Te�2\��W�*��l�D�T�(˕Z�Q�+k��[���-J��S٣�W*O+�)�T^V�P�Q���T>U>W�T�EĈx�$�
��Y"GL�E��#��B�TT�z�,�b�� n��V�M���^q@ϊ�K�UqL�+>�S�qV���Ʃ	j��_MS����Xu����T��r�J�Z��+�uV��X����������>�q��zD=����m�=����zZ=��Ә�k��CK�R�!�pm�6^���k���R[�-�j�Fͯ��n�n��Ҷhm��Nm��_;�=�=��R{Y{C{G��vR�T�\�R;�+z��'�}u���g�9�D}�^������R�Z�כ���Nߠ߮oҷ����.}�~@?�?����������?�?�O�_�guӡ:�	�dGG�c�#�1�1ّ��(v�;�W;<���*����gCg �Rr�b�z�ե&�]���
�����@��~�z�R���`V�_ ��$�23E֚��>�|Ch[*���G`U���D���h���=s����@�%8�p�y���/��`���a�?&:�	��e~�>��l�mg�OF0��ʸ�I'$׾�F/1[ �ڥ\�	���5te�x��v&9l�>��^G�מ-1���ܞ@��R��O%D���U�������\D�J�V˱�f���X������څ�B7����r������襬i�t�Z��\E��W���h{��0i'Q���gf��4.����|�,␠�P��2��+C�0�;ʰ+�?HsQj����)�lh����/N2���2��^�GIc?���B+�f��k�E�\�MX ����Q�A�k$5jo�/	����*��[ ��F����݀�Bu]�B��i���U������vD|-QXF��y���|����w�e��f@7a,��sG�G�[�iQ�+�������t�Mw��_��3�'4�d�K��.0�i]�k���#j������(��ZZ�����(��Y��%�O�`��U�i���J	?Kj�V�ה:�]�/ Hm��6���~������:C���T�`VJk���7�g�&1�bs*����^���R(�d�<Oa��(�$eW���?�GZ��ǩ��E���8����,1���1�gdY,`L5����Ğk�?��G�i����d߷#�W/�<���ǂ.�͎�.�ǹ.�Y1�`�����tD6����S�v�z�z�zbu��y3��V_�k��#0����7bJ�U��["ĺ�zK���mV�r7�W��9�8���8�t��?�_���(�J��Wq)J���LT�+��LY�,U��z�Y	*����&e��M١�R�*�Cʳ��Kʫ�1�]��#��rV1�*�D�H�E�&��X1Y䊙�X��*q����E�׋��Fq��Ol��b�x\G�Q��x[�'N�O�iqF�S�����CMQS�!�pu�:^��櫳��R]�.Wk�Fկ���ܪޥnQ��ԝ�u�zP}Z}N�����������������z^S�-^K��j.-C��r���t�@���i��Z�V�5kAm��A�]ۤmնi;�]�^�vH{V{A{I{U;���}�}��Ҿ��j���qz�������az�>V����3�b�\�ү�=�
�E_�_�߬o����ӷ���}���a��~T��������~B�D?����9�Cw��G�c�c�c�c�c�#�1�Q�t,q,w�:~���[w9�8�r�u�=4F�봻eY���9�5ᲲPT �&w����}��f �VWF���UV�jح��Bz��T�%G���������T�ٲ��X:"%~H�	���(�Br�װk(�.�ɾ�t]FD�e-C����Q�*!G�Pe�s�`�O���*�%_� ��Cfh5��ʋ]����z��T���)�@�_B%A���&�.�e�	�L����ms	VF��N&�Op9��UM��C^IN��y��V(��&㴫4y���d�m����4��7r�k8���Y���ˀk2���Q�]�)�Q1�!��}'�1�	�>|�*#�*�oS"�[�C����V�$^���/����ڟ�2B.U��&�L��i�P�R��]�����a�h�����S�9#�#FJ�nC��Q�U�6*�r�(�oW��1� .�����a�&m&^���N�	Z�Ԓ&�V�-w�O��I
}ɮ�K��l!�4��I[L�*w���IA�3A��}��x愜G~B�3?��:V�*�w��`�*�ګ�~i��<^��(<B�}Z���Һ��%FQ�t9�>�.�(Wy:8���k��7��OZ� ��eB��iq�]��O0[�}��e��⻒O�م��It눧��P>�����!�{گcv\����%''�>�^��ه��^��'5��J��?�͢�Vi�:b��&#�|ɏR��Hc�6�f�Gx�R�J[��:-S?�X��`M�s��q�<B-��H��o��o��,p�x���CR�B^w�G�!ʷм�EC$��%�$}�V%�~�;���Z�K���9u�Թ�&Q���4S���Q�R%Y*g_z6��.}�!]�}�N�1�r���A�O���ԗ)8�jq$�B�8������"��ƕF>[g"����O)���"�P_�^F� Q���*��	<�~�k��c�d��g�b^Ϋ����W���_�o����>��?�w�}�q~��G�o�k�m�����t�1f!�~+� 8��:�;n�jS�����o��"������<U��*G��N0'�m�n�.��oS&�����n�$hIji��o�gݷ��k��	�Dþ��,�j���^z
��ʵ �Gw' =��j�t����<*����� Wj����M#o2'���~�h#<���1��.c�_��q�wc��K��D����d���)�u�:��?��i�/�6��o,����X��32��3�1V �a��l�X+�e���>����αɱ�586;6������J��m�ٹǹ���{����Ϝ?c~��c,�<�|��:�r��V;��y���o��+����`��72��Y��J3�~�d��ۑ7!oe�~�x�.d�
^�����E~�%�W��6���89�_��$�C��{~�)��="�Xk��m�\; �^�s�� 9^e�ػ��;������c��o>T�D�e�M� ��s���zJ����(����ו�ǺT{�'�W��BO�=��q�{�ʱ�s�$&ʦ�mӜɿNFL�,�RmB�Jԗ<pqhq`�q�k�0���^��Yc=k�I���Yc5=kl�zj��Q���9��^�g��E�N�_�q�ȫt��2�Yyŀ����@V��*zYMO ��	d5=���'�U�'�<��L�<���q�l�����M�mhv���� ����5�j�B�K���V�-�Y�9%��YZ�гEI�hw�� �]�y��n�}-���r���֕/�_S�	߾���R�[��9��mz*�P�1�yB>MFy����� N�n��F�1ӘceF���Xb\mT�F���h4����Xg�`�l�n�e�kl5ڌ��c����k�3�;�9�p~������g�F���H1�����H5�Í4���j�u�����hy���$W �Pc�QbTU�Rc��1Z���Ƹ��`�jl46[���m�ƃ�.c�1�8�<�<���y�y���a1F��d0���22w+,F]�(��W�W�z�㌬���!��b��u�#|<�R��o?m>f�
c�q�q�Qc����ڸθѸŸø��l|���q��#�����P�Q�Wο:?v���w���0�=�!��1�H7F�C|p�J3�$-��9S�9T:l��� y�j�)�ų$�I�O ��N�����T�8�tP�K�K߄��g�J����d0a�����ǁ`5�&�!ۊ�yy����7_�L���	��!�
endstream
endobj
28 0 obj
<<
/Filter /FlateDecode
/Length 265
>>
stream
H�\��j�0�_E��Eq��@!JF!;�l��JjXl�8y��V�`[|�~!ɬ�^:�<�gD�F���ŬN 8)��~��[`A�o�ǹӣ�����w�����ItJOp�n���j�Ψ=��i@�
�r��g�d�N����1h�2�6��%>�m����B}
���N����T�(����<k�)n��e2�3QE�]�ș�D"���,�fI΂jVT� y����>b�q��%�չ0�y<��4>��U��
0 ���
endstream
endobj
29 0 obj
<<
/Filter /FlateDecode
/Length 1078
>>
stream
H��WMo�0��W�\��H}E�4K��v���z���a��d�����;�+Yq��'�|�pf���^f.���i��?���4��0;j)��y�i��	�i�k7#��[����O����$��f-��v����^(���p+��t�?�R{�PJch���h�_ѵ���u���=]8���CϪp7�6��|���&�=��*��ɋ�ެ��DT�t�{�` �zT(��'�\*F:]�l�ݵ)��N�]{A���_�>�m�!���a����Q{�����@'|$ ����,q�xx|M�6N�y�8y�kK�m���pSc8��t��~�y�j4��� �&�Ⱦ�����5]&Y���yL�U�٫[�މDn(���q?����?���P8��Q[r�N9g��B�� t�9rk��ܣ7����e�b��P&��;��ʽP-���se8C�P���<����	Dvw�z7��J��[�<! ���RИ�o�"`�(����l����x�n�
:B��jXEi�;dd�eƶL�AGiT��*�ШQ�Ra����T���*���OfeP��.��3R%��!��.g�H3�h]MAΡ!��˧��:F���TwQ!?����V�OE�zD���`ͳs
t���E������5����6M��s����Z�@��ΰ�YC[���p[T��Z]�>���N�i*Z>�Ǖ>'�2�/�J�G{��d�e��JI�3���@���18�E�R��M��Z��Y�/�����Mc��םb���`����"@�E�
x��,�^<�o�_lv(K���S[�TB;�S:!K˴�V�"����B]9�k����w�x�o�
�-��ujw�K����6>���-��
9CFML�9�wC�d�,G|h��5���̞5��]A]�dP��y"�}��#�G�#�(Y?#D9+�o���Ӂ���c	�: �K���>R�u ��z[��zU[���R��M���ʓ�"�k��Q*�m@�􊤬�{8M+�����f\�;�����.Չ���]7����1�ɒAͳ��v�0 "��
endstream
endobj
30 0 obj
<<
/Filter /FlateDecode
/Length 772
>>
stream
H��WMo�0��W�\��DQ� M�v��0�0�������H�Ie�igY�6��Ъ+>Q���n5~}k�G�уq����zhd��t*��s��E��N������ȟ�F��q����]�Jo�6o����۾t�o�,�k�C�V)ev���_�QQ��C�,O�:��IR\h�pu��.ާs\�].�Ac�����&�ydq#�5�u��Ibw���X[~0z�����EXȸ�n���  ��	���`��E���H�A�9���@;�q�.���J�O��������� Wt��A˯C��) Mi~Wr+�t�9�ɋaFc�\!#�P�.+�m�^����9�.�tS\+<�U2`�A7%D=��ե;����ns���Wܝ\R�]7�Ԓ���"3�kf�j���eR�VM/����	d��eE0���
D'�a�fۿ?Ô��Y2Ǭ��P�e*`#aN�e�8��T�.#�Jo����g�A��ܗn�s7��x��Ҩ��m|5T��6VFm,;ǅF�`�U��'%�CR��QlJx�m ?�]A�u�ik�� ;�q�`�%�	:�":fkE�Sa�Q�CY��*�v��&�tW[�o�D�..#��U2�l����Z£�d�ԡWv7���
i(
��ʱ��L�r�X�O �tQ�hi�D{i�$��Ő�%�h���䭲�z�5=#�c�����ȡe�%k�L2i����PQ�=��򢛜=5�#��<|��(\�<��n�+�fw	r����-� ��yy
endstream
endobj
31 0 obj
<<
/Filter /FlateDecode
/Length 809
>>
stream
H��WMk1���s!�f���顷��J顐���茼�Wڵ�%�氘Ĳ��<���=���S�Bo�^�c���
���}���N;!5�����L=�~w��7zm�N
g���Q�{����þ��IJ��;/���?)��dCk�t��7?����н�z7�\��`~�-G����`|����V
��D�6ß�-ΐ�#���2��$zl��WS��nJ�-b3�eOx-���E�"��0W�"��V����J@Q�h�j���J$=a���A+��csR{�lqUR� �@��O�iE#���7a�&>�0�(�J̳p��,�(��`�\ RR�@%F����,*y
Rƙ�m�Z��[_,���pm�4(|�-մTCYI7i�z���Fi$�&x��
��:E��8\��h-�k��k��+�uU��H�XT��,�����␕�Qyw3�}��@��-��$o��V�YK��\�i�V� �7��}dc����^��#��eTN@U��0]��)���q��lh�M>"�TP�$������E�Ǒ5i=?(x���ß�D Ys�+�ܦ��8G��$����t�>��t�ԥT�2�	����%�4/�P�E �,/ojbgT�Kl�����F�Où�=�� S�tX&���dq�7U�3h�o�j=����pk�5�{	w�z��m��h���#����U�#�Zm?�$���*���<�������iP���!�7!	�����'�m6$)�*�!maD���.q	��E����T�gX������  78}�
endstream
endobj
32 0 obj
<<
/Filter /FlateDecode
/Length 741
>>
stream
H��WM��0��W�\ة>F�ئ顷�o��Pؖ�����ٛ�R�ԒRv�����=�h�̌����=v��]w���?v���Ϗ�>�{zT�핳�����n@��߳%�'q�~vo��tmp����j���/�
P�q,��{'�л��j�UJbƍ؉�d]�v���9s�B���yB�� q�u\_�v UFՁ��4k������"'"x��N�mB�kp*��G�Բ̛t�l�5�;��;�8���NE�N��,ɷ{��3���!᪄��\z��g�8!�E���H_�x��8(h�����oP~_q�}�Jb#%��h�����Lu��h�Hi[�zr�	��m�`�ʪ�8��a*�K�EvÜ�Ts�䊲�'4o�6lp�����k��Io����[y�?�"13�/c6p�Ԏ��<1,���T�0S���d��(�:�{�����>�ퟝ?�y�H)��?~�G�ƴ:��`</�6������*�I�Y4��yP9���@y��Xf���F�҆�\�Zp�)������xqD�5#RJ��N����g�i���ANy5���ᘸ},�2Hx�;���nP$eH����[FqM���Y�0��Ց���e\}�`
[��պA4�F+�IQI˂d��O%�tM�YQ{�$r�R��(�@ťB[�|o���Z�@^��}U�(�Y>�V���1)��3�������� nz�
endstream
endobj
33 0 obj
<<
/Filter /FlateDecode
/Length 898
>>
stream
H��WMk1�ϯ�9c���@w�z+��ThKi��?T���Lڬ쥇�e��=?�ѓ�2�nqY[Z�\�A�1������#}'ڤm���bt���L�6)��V��Oo�As��1��&��m�q4����Ӈ����?=��a�U_�P�F������sA�ߘr�R9Ǻ�=�U}�s~h}�j����?@yV����O|(<��ü�D��7lG�<d��A3��D� ����ma:��"���k���X^!�h/��.̠�� �CwU|R��@���6���3�J��c��^��砭~�d͛*k����4�,��z�iuY��|)��»w�YǶ����Y�V��+���:n�)�ѣvv�8-8�v�6�~S��+�w5���u�壌\D�S�!W�7S��8�eoI�cj}��)P-b�]Dl����Z�_}m=��M�a���n�b�Y�93_3�Zԩ/Y�N��M(�B��ķ@�!�ɷ��|;zSv|^�-��U�{2��[�F����?6:Z�������*=�Eh�egf�#��eۢ(����l�}_$TaL{}�Hr�7}�t�'c&��5n^�	:D�w�$q���"D>�<`�}f��z�P&"K�A�"d���D�9��Ȏ`&���-�NF�/v>�B�a싌i��VFa�{-신^=��f�M�*�
����g�<�>�
v�_/f@D��zP�#���t���X.�sS=�m�]�tn�	�.�<�B-�4��Zc�Ö�-���?�)"F�-�� �-XWP6DR��[q�##`h���X��Y��?	�n@�K���6ʠ�$�$�G6�@�jri�0�DD�ny�	?�"�����Q$�'f�e]����iŶ�$m���*��  �M~�
endstream
endobj
34 0 obj
<<
/Filter /FlateDecode
/Length 949
>>
stream
H��WM��0��W����f�i(�M�z+䶔
�R����?T#9�$�)�xK)�1�e'��f����{)�as���.�&�0&lh�曻����n�^:)��e8�Ǖ����AOǯo�K���p;8j �5�C�ϝ�;��L0B�p#ϫ��S�)�c���?=[��^h�k�`|�F�6�7CDi���
��cZ]Yb3Z(̰=F�s�=��F�����["w���obUk1LYmG�p���
?�J����1	31�a+����ƶ{��S�'J'p�D"w��_�YL��:�.��	h}4�V7�ŔE"ot��M�Бd�0�2
�)抂��b���1�*��y�qAN�BKx�����^$���iy:Ա<�*�Ѩ\���J�a�`N�C����GS(�0���k��$|�*2��⊠b�+S �����&FU` ���uU26�MUA��j�������ۤ��_6GG�H�_��Uf��� )�lakS�h,5v��De�Ʉ��<�ur,�L��L��k}���U#�q�CZ����SV�т���C��<�U!���T�l��d#s�CCe�m�y�(��Γ|"��rsk>h�pu��٧Yq�_^׬��{�a^q���H�CjԘ��=/�!��n�qbI�х>��@
m���4m��4O��y�Dqav��l�䛣r������A%������%*�i�<G_1؁b��U��T���F1`)�r%X�OA8PaY;YP!�F *G���(����*�w;�B/���ǧ	�����B�B�-�� ��@B�o>T�X��c%]L�FGЗ��/� S.��9��*Ɇ�R�#f>����Tf��8.�}�����Av�Z��7so��Ws�-�9i�]�zbrj�
A){+��*���*'��a�8�5Y�\2�,���V���n���~�u���` �w��
endstream
endobj
35 0 obj
<<
/Filter /FlateDecode
/Length 744
>>
stream
H��M��0���:VՌ>%Ф�Coߖ�Ca[�������q#��v#)ݲc�X����h���;�������2>�a�Ώ4����t��n�e����c���B�qs�ŷ}��_߻G��<��tA��2������ ,O>��<���w�����~�	��vb�?���/=�aߑT��?/WJ�-.�j���N��Z��bsqN:��S�eĭ���띰
�
�P�t����i3p�i�d⧹D	d���p�q��hw¶hwz6v�����Z9��[ý�p�\�C�i��?�U5,&`PZ�S�����r;Υ^��3��H�����D-k�� zj��)�g��IC���K\.�%^�OZ
� {�"3Q{	���8�F���|g������/ϳ��<�M��gs�-x�>q�ŭ�Єq#^�g�0u<�{+����]�.ܸ.5���p�-�9�=n�j��ĕC�D��2�+S�%M6T�S&�
�� ֙2��hX�4*�׉��j�cxҁN_���� �A:��Kl�����fo�i��O׆gQl�ũ��k���
S��&�@'�RZZ�S,*�n*�7�EU�o��5�C��Y�J��-�A;.<��@;�Y�(��騳�-��L�u5i�
�ɬ4!��0��";m`���L������X��9�jCð�:jU�(q�ݖ9z`�V	:3fl$U�
�̔���2�q��5ؿ���x��oIi�ʎ�Q����f���W���[� �lw�
endstream
endobj
36 0 obj
<<
/Filter /FlateDecode
/Length 942
>>
stream
H��WMk1���s!B���b�z�Vz*��4���:�];�VIXIΩ�Z��z�f�|<Nϓ�̒^7����?Mj��ߟ�3}�}5;���=e�������S"]�����cz����rT\8��UB�|z��~�R��/�{�s���e�?탨�	��S����mhQR	L�!.��=��Oj>��P�۲z�c��oK�N�/܇����H��z�K7}�q����쩦P 턂��Nx���Ż�ˊ�.�t�� QTD�-_2�e�CT�k����3w)���N4'�Pu(���Z+���L@?F$Z��H����H��V$�+0�qI��`-?:�V�f��Z����;%�&�e��7��tF�p\x��� 2h6�*��@,��1e�6��2��X�Pͅg��w7N.���Qv�����>����H~�ڟ��ƹa*`R^�B\�D3�)�){���q7���`�p^ݟ�1��_;V{�lݱ�˱����󂳽ֆ;�Q���<�e�=�y���]y�ۇķ �|k|l8�q�b�5¹Ա�^��� c���iUT��Dk�8�e��Hi�ʨ�kg����D)}=����k+a��B��<�UG}� �����6�b-m0�����Ыځ�pVmF��"{T��fU�)���[H�g����(b<��z�$�3+�|7Z���6���FD*�, ��ό�)��QY����br`ZLC��!��iߕ,xo&=�ų�i����Ai��8�S�2���r�2�Y��`��͐��qc�]�iǠ�LC��M�Rx���W�Q�S6ך4z��y\V����>eA�N��:4�+C���pu&�c:���V�:ǮS��׉��䐋!�6\cK�(��=bP��~A���k�-�=YqiVrF��b4L�6]�;�(fy��!����& ˖M]���:�` !9m�
endstream
endobj
3 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 4 0 R
/C2_0 13 0 R
/C2_1 21 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents [29 0 R 30 0 R 31 0 R 32 0 R 33 0 R 34 0 R 35 0 R 36 0 R]
/Parent 2 0 R
>>
endobj
37 0 obj
<<
/Dest [3 0 R /Fit]
/Title (b764a1e1ed943a36a59006d6520736c8353323b5acdb0bb64bc57c36469333d2.pdf)
/Count 1
/First 38 0 R
/Last 38 0 R
/Parent 41 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [3 0 R]
/Count 1
>>
endobj
41 0 obj
<<
/Count 2
/First 37 0 R
/Last 37 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/Outlines 41 0 R
>>
endobj
40 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227170530Z)
>>
endobj
8 0 obj
<<
/Type /ObjStm
/N 19
/First 141
/Filter /FlateDecode
/Length 3662
>>
stream
x�Ś[oǕ���+��F ��^��86f�	"M����($Q�h`�ﳾ��X�-H���<����ڷ*�m����ַR�ֶ�Zݪ^=oI�ږT<�����
�Ի�x�-�m�>���1����em��]ǖ��]��H[N�X�lj2�k�Yۺ���/.��ͳ�7���o_|��������_^\�������7?o_|����7*y����/n^�Ŷ_|���~��G��\�����'7�[ڵ�?����w7���z������7��Q����/���ݺ��W��|s�?��Q^�k��Y�*���~y�B����ۻW����}yTܾ�)[J1%��~y�]>y�O���W�^�i/?��~m�ܿ��������޼�~�?�J뮵}���ǯ_=q��^>��y��m�z��k�Ns6��������ӱ�Zƙ+�\�����[
��������_�{x����ޟDpq����|�5�3-X�{뺸�a;�۩���4����չr��1-�r��%�R;\<�]�&=�V���d<џ1�+��4-��2�6Z��J*Z{B��Ҧ�C�]˩i+�(�(T�Q�^��u�B��Z�4A���˶�.=�R���v�Ļi�ز�Ho�� y˼�֪ճ��(�6WU���)�j�-F4�o�D�\E�Sv�]���Oqp�MJ�1aL)~�i���C�5��ؓںB��K.L{�ǈ����j]+������D`-�+la�R�7��AS}��2���b��-��$1�2�l�i�NL&dGm���h�p� W�vEC5�[SH7Ů��������}��B�G_曻�ƞ�R�_7L�8q�� �E��`ISVp��i�*��)*��Fض��$ I��i�$�/�\mXh�"˞�jN�Jx���.��IhP��w�"k3'�A�bc�
�����*��	pE�d�s��Nl|�kf;ֹ�;�E�0�q�P��j�Y�l�����ނB�gr@I3hCSlȝ5��`��!1O!hJ���u��3Ɨ,C4�!e!�0�!�Rp� kg�6ش���	�X{(EF,x+�1�&#����&�_'P�.�1!K����<ÐjVn��j��R+0���T���[��<���V�FyC��(ܨ� ��#��ZY�V��D\�1L#�b��h�G�T����%�yͳ��%�#ڻ/f\
l%T�!(,�B���vƙ6�F ~��I�wE"�ޭ
��',A������
��jP+K-k�V��5鷭�-����	���0���dUȸ�P���S�Vq�j�,N��ic%Zh��b��8j�/�W(pߎ�8F����bGԴs߁4F�0�]�|�K+�+}a40�/BXg�D�L��]I��.}�k3Q��*�qG�'�����GC�1��?�nS���R4�5-h���0���}���|m�y�~���Ց��l�^���S�yU❈UODv4e��BI�Dy�ͱ�t���c��U?��>����*@[22�t�fpl��?h���#qNF�*��&��n
+��-K�8��I���6L��k��#8�җFðZ`��x��C�41K'Z�����U�-�^,�����{�ɘ��M��u��t̼e��v�׆���꩷� ���ˑ�$܏�wI�$'���M³��TuX{�@�,Ç0�K���6;���٧UJն�%�(8���t�T�$�������k��<0�,�?"����}�T�п�nc���U,ƨ��]ؠ �w�#ֱ�k]�Wa��5�Ɓ�'t�	"���N���ly���Ŕx�F�L�t���!���6���R��z�6�m��;�"c<_ݣ�(W�R����=��d�T�@~�q��N�.�/�h�\DB�D	Q��j��'-��G
?:AM�j$�q(� �ǫN����+f����μ	"����OL�ȁ}t�ֱ"�&ܘ�-Fڱ��M��K������X��wO):xf�B��g��g����آ���@���� ���"k�(��9#�j�f#<[.,��G��&�0�0�Nvq�Se�2��پ�6�.�G�MSr���Ϧ4b�xNҤH�����䅯=ڮ�;�>���b2��iY��[���z�Ζ �j�~�J�9�¾7����86`�˰:ҷ)m\h-�vw?3zf�����/�#bP��͞�7�bW��f��Ƥ.�x����.�u�_d��3?A�ȶu����o���`�����wq��!�d�kG��c}�x�X��XC8`��;��2E�]5q �#Wp͙%W�L-�`��`�^�9:?#�#�wTc��{C"�Y�c���r?f 	�q���\[���1�վ�3����z��D���^SJǪ����F�e��G�B?$햤pI��I,�O���(1<N,ؗ`Q�͸��������Ev�Kd�Ή�4�4XIyTL~��q���'�<0G����T�ib�g��Eg��q!w��j�'Y� ��H�%����&���ˠ%��/�5G�D(���0T��q�1�$ �X�=&�����RF�d;�D�JhhK88)G6K�D1�u��0ϸp������G$�$�f�K�2=�J'U2oV{	
�����������i��(v���(���n.�2E���P�Pm8�<��g��]?��3)�8o+2j-�s�X�46E�� ��B�
�%G%Q��w����QԽ8~���qq�B����#�A���[qj� ��%iZ�i���3����f���K�:vd�����;j�q
G������`�4��H�["��Ӵ��#q��y\1�������~�oO>w
p>��Q�0&���+��D�l�|\��[jG������?&����+�%R�D�f�;Ys,��<�9\�&��'�C2�q�|�C��s�_¿�R�E0��Af�A��q����-fD|�Y���[M� G\X��"K�_FA�y�x����D$~�%��ω$��"�OGO6��Y�U���$oJ(���an��m���lb>�9O� ���f���%�8�۽� ��b���3�#�u� -��qj��qbӏS�F{��+.N�C���B!.X�]����ۭŝ�������;��˝G�=�I8_!����[5����~.��7C����#��#�� �p}!��$;��Aᵃ�c���.w�wAS�w^�8����L�1�9kPD0A5S���;1S����q
@^T�1��sAuSc+1��y9�8�7�a��ߎ�S���
E�`��őMP���4��xD?Pݏ�b?Pˏ��%*��c��6(�H�"���\S��&�[P~L��j<�:�)2��&���c|�<��t���PK���_}�>֋�盾'��ը���k���wr�ߊ2�ӻ�|���ׯ���G7z/O�|�t���R�Oݖ���ғkPk�נw��;M9�T���&[��}c��1���W_]���&����y�OB�l?�w�����T��!��.�r� R�_�����CH��YH��@*��H��/@�#P�o�l���{z'N(B���o�����g�pG��{m�����������������r^��� ")�
endstream
endobj
42 0 obj
<<
/Size 43
/Root 1 0 R
/Info 40 0 R
/ID [<5217C64AF857029729064CF134102380> <A09F69FFD4BE88859A2E12BF358F174A>]
/Type /XRef
/W [1 2 2]
/Filter /FlateDecode
/Index [0 43]
/Length 150
>>
stream
x�%�;
�`���GbԨ�������D�/�1�A!�E@�o�!��X���`w���b�|܌����&b	0��ȭ��H_�k��h�&���H��z��h��g�"�NK�v���q�1�~�eb��6ʱ���@�6�}���z��
endstream
endobj
startxref
54389
%%EOF
