%PDF-1.7
%����
12 0 obj
<<
/Filter /FlateDecode
/Length 20
>>
stream
H�j````b>�	  o%
endstream
endobj
13 0 obj
<<
/Filter /FlateDecode
/Length 1201
/Subtype /CIDFontType0C
>>
stream
H�|�Lg��Zګ������i`�2D ��D�8I;�Dc��Qۣ���V�jJ��	E
�LQ�E��4�ը�?�"l�G�E�Ib��{��k�ϒ%{����<��~�<O޼(#CP}��|����,Vo-���8s��I�����U�b*Ίi5���D���m�'�9bB���Lq�:%1�:QH��� oP5����o�t&�j��K�
�`1��ٌ���ԈfD53��0�٩lfzzzT3�:��z�z���m��:��*x�`�Li�-[ب��8'TE����Zl,g��qk��f�t_�L�]0���a3�G2����)�Z����[-�ۥ��5XM�$>Z��WZ킅�����9*86�5q���4��H�"��K(-��Lp%r	բ��92��|a�wD�}�4yD.zޚ*{�*���)�������_!";�p�@�`��ENJ���ѳ(���q/��%+6�nٛE�S�.w��� {07y,�����D��k.����B���db���� }���w��rZ�aƿ�L&��,��y�Gњ��'�� 8���� �)X߇W����5n��Vm��]���e_�ogw�E��{~��4��"�R[[�ʠ�j����Oя����Uu0���J���7�s���12�J�����O��}�r���x/Va�S]�gT�"�]��:8.) '6�+wn���Ày�z����?ɸ�>��j���n��kۘ@My�H�V�KmI�6�d����w.�.К�-�B�y72��8��W��v��A��2��QQ�T�B�Xi�vgI�ʆݯ�yt$�gcx��nm�E�D��(d �:o��x�WC̍��c�C�=M*<�]'6s��Z�� ����๚����3���s n k��Ÿ?���1R�]��m3[5�7�Z�����%��6ћ���Pq�]w���[4\Ɖ�gז40��n�oeQ�������aJs�yFdΠ/@�9���D:L��@��P�&��Q�f�M�̞r���T8&}�� �h�ŷ7o2���Z���:��~��o (��j�s�KU�}���ՑЈ���nz�ы�6�7�&�>���s�d/u�ݽ���o4���>����<j뵬ݨ_���D���"�~g(1f2~g��;��R��6%l=����{7��yձ����N�D��[� �K*�
endstream
endobj
14 0 obj
<<
/Filter /FlateDecode
/Length 263
>>
stream
H�\�ϊ� ��>��C1M��KK!���f��N�B�b�!o�-]XA��|��7��^[��oe�m���.^"�8jÎ9(-Ã�)'�'s������5�O*����{Q��=��^��f��������8�	�AӀz�ML<�����<���!䑏�i�NH���V��V�Ш�sr���~S�%���(�HU�2]nT�%e��ERVIYf�n�N��y�������A��=e�s��X��s��: ׶ٯ  ���
endstream
endobj
19 0 obj
<<
/Filter /FlateDecode
/Length 22718
/Length1 49828
/Type /Stream
>>
stream
x��	|TE�7\˽��$� lI����$�Q��!` ,!	f�,l�l"[d���Ã�0�0F@@Ee��]G��ã�&����N:����~���?�P�֭[u�lu�Tw�&� �grr�芗�]%��J�v�����݊2B��q���1�΋���(!����0e���	y� \�������Ϡ���������"B��ٕ�+�M���!,&�lf�dv�'���@��3�1�	@���g�˟�D�B����Ԃ��\���?����h0�2�����RP\97ő�@��g��d��_�%d���g�-�e���|Β����DȌ��]VZQ�ZB&��S�<�l�+'@߹�S�+6��fE~�4�!ߓ����s������T=f�[�xa��X����jW�zLR�~)�ŧ7�!\�3� [u�4���z�������ƕ�G�Y �47+�)#��ɿ~����c�rIq�\Z�H�����	������-R�����ُ��ds�=t
�M���K��|��\'[�*�֡��ZD��$K�5ҁ����8CD�U�UR���*�Va�M6�� ��N�$�t�ڂ�K�y pJ��0�#5�r
t��Ut��yOa�Tp�:���{<[C�L���

��d�G_z7�ZM�`�,�
�_�^/M@@�^u�Y���M����p<=
ޛ��[
ܰJ���,h�
 Y�,o,k��]V����mJ~�"��$<hY\.W=ty}� g������:4�=kd;YW5�ė���Q����o*Ѱ�����+�.���y�)p�y	�`h!S!�t~KVJ�YE��W_ґ�K{�H��y:I.5�$��i��u���dv#?ҕ�$ۈ?��hXH~דd!�t�ŸԿЗ��v��o�B�[�u���ֻ�E3���9���U<�V��Q�,m.$��E7`�=	b��UD�!�0�0�+uMZc%_Ĩ�k�5ך<<@N@ϵn�&���� 4>�ç�w>B^�,�� � f��d=fM"{�� ��,p_�o�aQΧ�f#�J>t�4��j�4���z�a�~O�dk'�����[ɟ�
�%� 6]�y��x��t+�^���:�&�*�0Нvg]�ݢ�y�C ����F3J��]4�f�O�p�'� ��� y���m��B�F�#�b��4tC�x�6�\��Ĝ���s����Ig��4ԯ�Cr�Z��fxG��ɱ�2^Yd-p41c�8�c���T�+r})|�K[�"�c�����
���
q�I/s�A�˸������W�G����J�����EUX�������>�m��Y���"֠��$�VIv�u,֓�@;�3�L�=��Ur�&�
��H(�� �N1���?!��C�h��N���[��q��1"���u���]� �h�
�$��|���O�
���H'��� �����	�;#�H*V�B����]Bj@|�n)�)��g���P_*�����3r��a�)��rO��zh�����-�x}�A.q��LB�"6���7�*�A4f
'Sd	�|�h{�ݻNr��J�c����x�w�[�"B��<5��(����ge�C�������IO�m@l�m�M�u<J�t�L���Yg�q�W��}@o8Vֻt>��΃n�":<OR`�]�o����Q:\���H~�g;HV@���[�x��"bCz����	�ݍ��.�޽��*�E�.�DPB_$�(�1�c�$w���u��p9`)��H�:�!��L�����ch��Q��`��.`
V�&��aX�5\�$gi��fM�c�,9�!9]����^jv��%��"29��M*`��a�Yd���9�<�Or�>+��~8�����/���$�U�M�)�����<�q��>龊�C�ށ�q�� {<��O������v�����h/!54�>�{v��=V�K��ԓ�� @* ��U�"�&�t 
Qϟ2O.�-	������)t "�d��B���t2q�-��@��L��t0bY�e!�Ƹ	����l����>�Q�6TҚL����<u"��Gϩ����Zم�x�*OY�zgVW�ǓQyJ ��J���k����R�mqci��1�,F6%�ݲ�T6u��j<e�̄o}��"����Yb?.��xg����S�s�Yy1�ȧ����%� �֋�"W����k��5��Z�Z԰�a�nn�֘��5�5�!��a����`��G~�=�J[a�cw5�c�}�>��z��57�'�ՈR�@��IzPK>1&_�y^�/�_��,�H�_ #�/)���^�/�������Qw�@�
��d��; }m}-����?���M���_���~��'�Y���Up=9�"���W��n��]o���8�y[ù�6���Vfap�{���Au(vS��^چ,v�It9��qŨI�U:��uyRA����]��%��G�q����$D���D��s �y8�"b�FT~ ;�8�Q����{G!����/3	+�}5|}0����pv'�܋�cs���zKK��Xjݐ �h|&��{����Fܽ�V���)kc��u8�=���o��<��'^�DK;��w� A�qߵ�*{�"2�C2'Jq�t�$K K���<����ݴ'<�.	���`��)}��@�~8�_gA�<;�O��f����ϓn1�nii��w��2��>0�놖#;ʱ��
2�,���4��|d�2��~�̥�X+��p�#
zf�O5��n2�dA�EaYF��g4���(���@���zZý�6�3(H��h�:�N�v-��v�&j�k�Q�.ے��pϕ�6�Ў]���� �=���3;���P(<N#���ձ z���+��ύ>������x�p�ѹ�Υs=�޾~+� 7~Z��@�A�I�]~X�o]uJ���~"��n �u�	�lk��T����R�D��]挀fχ���i��l��ϡ
�E��<��ED�sQ ��(�gf��9�=��8�D<�@���.���p������e&�t@�r7�9���Q@k��}8=�"�B��S�ݠ9��Ӊ�ð^�p�X�q���F�9h����bq2��ڛD�r썳�?���c:�����©�N	����Bf���xA���pV�S���Z�6������(��տ'��`����n2����rZ�`���!��=���z\��nG�ն�m8Nb�P�P�F��lЧ�Ǣ_{�b � ���6�p<q������<uAT�ڊ!=Y�g���w�CK.D�(D�xйJ��|Z�L?���3y��
h��a����bpy&�.���I:X������w��E��`����9��,�	 g�N�ч��"3rm �Z�]�JF��ж�f�s�����x�:�v<�ϒ'�T�9����������8�F�,d�L�M ��w �a�X��@���o><�K잫`�0�[��+��C�Y�Wy���+θ�E!V�2���w]4"�;�s-�+>Q*���%e<�8��Gz:�D�V�q�����~L�������+<|����K�<W�~����-��u>��}m�K���jv=%�� ��.%�=�{x�W�#d�����#�O���?�L��JG��|j�}Rr��o>@&�N
�dd� ޝd�f�#X�wc��8Cuskx�?\���]B�����:�|�p��짢�O�"eN�i�0��T�sw�>	"�5�U|2��X��c)$E���h��˅��O7ăa�3��'}JH9�P������I�g�|*w��]���2~�̇8�F�_�9ŧo�Ql(�P�q�����2�]bPƠ�sR��	��#�b��E��QP�Q�>��R�.�F	Jʽ(�(�P�Aǽ��]��I����a��R��HO�Ǩ��~A'�H���u%���϶B�j�}�-v�v�1: �v�~�un�����[�Kh';����f}�F��طF`g�=4U>:��� BF�?�s2�B�/y�>�}�ot�<o�T�#��t:�����q�f9�N��+�ŭ�ar�'c���sֺ\c�����j��<ܼ_	��~�+r��,g-m���&�4=�Y��;4�=)Q>��W��/e�~gN�s�cu��Վ���^`�i��S�;��؄9�b��@���J� 8����؏l��u��ƇS$��>9���8�Jz�ˌ$�S��k��*�l粅�7Q���z�����_G��������:��r�����j~}���������8�Z���h�����h�?:�����o�?6�:�X��Z�[q.�����Wrկ7�+��+������t�e�W�_����Ϗ��>m�~v�ڎ����t����u�Ak~i����տ����6����������"n.�t���V���m�o�����\�ّ�ц�Y��6��ׄ����5�������+:Y�g����u~J�'u���O�މ@~�Ώ�xD=���ާ�x���X9z$\=z?�	�u��&^�.^}^�p9t��	������@.��/�����>=���^�{u�� �G��>�>˟��O��W���w�����K��|W/�_:ߩ�t^���Z��w<�Pw��O:�o�|�Ο�$O�|�ߺ%Jݪ�-Q|3�߼�oz���I�÷?�_�l\�n��o�S6��1�?��G����|��.�?i	�km�չ|��&����t�R�+t��r�a�/���|�Η�'�K3��/��=�P]����|�����u>G�u^UiW��xU-%q��J;�<�T��8�\��y��KK2��M����Z�����"���g�0���3��|���<W�93���� uF0���t�O���I6u�/�/�O9�'�fr �d���@>A��u>�C;u\,��y���u~�B>V�cy��G�^�h��᣺�)A��<eX���G$�#t>w�sy2� ����|X��:,��eqq%!�OM��	���.>�W���������8_WK�n�ݢ��4..W�G�w���o�!:����AP�\>�w{u�(>@��{��u�o��^�;������c�1V��w{ӞG�ģ,mԨ#�Wd+�W �U�Ĵ�5���nRz�W{�z����`��λ鼫�#�xx�5<�w��a:��SCu���K�;{�Q<3뼓�;B�u�V�Ў��y;��-(�M�mZ�R�$�ց�u/��ЯU �� ��Cr����0t��kW�����;_��k羆�|�;+���*v����tn�$V�[�p���t����s5�s�obs襲���ڋ��4w�Z��������!���E�C�5���lr6��xWѯ��NW�è�&���ȷ��_A޿'�Jg��C�/F��#U�(y�P��1��C:�O@mU�,\|V
�~�g�4QLv�}�� �,%��,��,�����d)E]p��D�Lr�laW���y��ѱ��9�Ed���v7˗3�[�6���
�`+��g�E�TBBf���Eu���իxBH'�V4�A
����(����;T|B�ɧ����r%L�ï�u���8ſ�^��:SY���y�t	��e:�C���~����`�	9���452�˿9x��5�3�	�?�t:BI�C��E�W�#�B3���~���<��5���R��M�/�A�0��X>]n�C��<����o�rz|�BR��|(r�}�R��B�n"!GeEp<D��2�բO_��M�.�Ŵ����ٿs�B�+x����L�7�-�d��h:�á[I�B8]���f�0MQ� �tmH]l����{k�z�v�P�G��Wić���i���>&�4d���:�A�@��.�j�u`@۰֯o� ^�|ٲ�5�7nܬ\������/���>�����)���C�$蚨�L�� ����6���&�u 3���ח�)�f�ku��O>Ӈ�}E_��2}g�K?��ld�?Dj�B��pZj,�vnݙ�2K�l�.��%��.��Cd'��D_�$ZL�F�������D���]	� �ˠ8#+LX0W�%�Oc���s\���b�\��BI�_�p�
�ָ���-��훃6o��:��֙t�������P�|���ĽM�i?�G+�j�m�6G[��Ѷ�d(ʆ��Pu�6�4�<�2�:�6���c���42�NcӬ�l;�����;��m�i�y�e�u��9�}�=ǟS�S�Ӟ3=g~���9�qr�g��q�z\;n:n>n9n=nK�)f�S�i�4u�6�4�<�"&�)B]��Ѿ��Ķi���F�
e���>���U�0�B����1��Z�v͚���Y��?������v�}3`���R�v������~����t �����K���\��>Hɿ$�X�DI��$".�oV�fu��l��ô`��`��������¢R������K�����h���{���ڑ7/�!����};�{㺓�᪦�k��v�45�������M
�̈�ʨ5�m��w���\'N�rOx�\�]&�����ĥm���p�ݯ?p��7",T3�����U�3�/�Ul_}��/7y���g�f����M�xqϞ=gh�=�7�Y�H°s�c��8�De���j�
�8 �v#��o�ͭ�k,�}6k!k��;nۤmm�l�6�l��!�����_�s��:��p���8�C�i�@V��/���=i?�Ҍinް]���3ߝ����lٶm��G�x�`ދ)�����t}��7����~}7�]�u����u;�t~�v�x&�O�vd�	q!ԇ��}��6����P��������Q_a��#P�eQd�YyJ~ub��v�}�����s?��ޝ����W^y�a�ک�����}v��i�q��u�]/�݉���:��l�_�x$p��LV�l5�	���m0��GH�0�i�z��֗~��]��VH�@�LqB_o�k�{N���:�/~�s&m����t��{����:��o��ӯ:���ǵ�ph�g�Hpf
i����a���m�es�M����$�'Ԥu��B�E���\gD��W��{���b�	E�sb)�αmh��:���(�d�#�O�����\�H����������lܸ��+Ճ�û��˽_��o�봊>J�ӵ!E�w�:�����/���S�T��k��3�x��*	*4�U�i(	1���r3��V�Y(�L�.1u�5|o���0sC?����KԞ�ݮe�I���a$�����]����6 �v}6&�ޥGp�.�~���By�_���N�Mh����nt㥂�(,Kw3��@���t�1Y���/_��q��%�~{��o]�i��_���v�^<o��E�[��l^�z���U[2;\t୷,:ع���]��՚W錹>8w��%��/�L�R�.䮸�V���w�5�G�C��7�no�qj	�G�f�\K{6�����!����+쎍��3@X<4�e.ٰ�\���ha��>�ʷ�G��S6�MS6���ig�.�~j��?Ԣ��K�zE��A��t�9H�8���Uvj*�� X�"^36\��[_�t���ɭ46蟱oAC%�ʼS��Evj{�\!����fE� 8'����֚������3�r|��G��/���+�[����Ze�2��9.@U%*ߧ��D�tN+����kM�Qe^�>���'Jg��~B?�<ݹ��vɢӕy|�[F�R��bV�!����|M�}��̏�0�^�����rFTe��Ic�"�R��O�~T0$��t��!}�n}���n���#��#�HT\�v$�l�>�pl�l�[۷����ZL{!_��gĄ���X�m�a@���(�G���Ci��;G��3����g��M�׽;�D�h	�ڽ��w�a;����~>�n鯫��ӱ��ğt�k�m��$��4�g1�X{oS�#& �ԋR.p��������a��$7ݩ?=H\���"�s�x�����o������~�q��o�c�\���=����5�=��&�z����?X�j�mB��c�cO�I��"�>�!�=�PΎ��17yO�����d���t�k妭�����Z�dî�҆),����{Hz�Ao����H3	�{+e��M��'fN�T��}ժiJ�U#1>���~�t5w`|���<;�?+%��uQ�VK[�ۚ�,�;�0w���q��y�����r�e�:cK�2DP��̇!�ѯoտ?�S��ݸ�S�Z����_`�*��O~�ʲُon��ok����b�IF=�'�zr;�V^u�jŶ�+Vlݶ���P��
M���/���Z�Kڎ�������V�t��X���u���V�g\��@R�2�a5㠤���'��>��,nu�����txg��(=!.]�u�o���S������~M�nxs���v��G�7<c��u�ba�V��f���Mܪ�s����4���J��$+m���Ƣq+�'}��]���;�l��d��`��D���A��9_�NE�նU���Wɶ�(��V���_�~ ��i�u�=�p��Gټ��X�[/�󞺯a�z��7a�Y��U� �rL����FY­6�9�d���Ōd�$�X�%�p�Tq��Fl4�[�ͬ2�i�lf��T�ܥE���1X`��/7�g[/i�����=�u �:�GUlAjWڍwW#lY��l�:�f�1���́���3W{��m��86ќe�c�!����_���A�H��O?����^u�^����iH��5,�m�gcz'�-]����Dj�Y�9�i	��֏�z�ر��E��< b)��a5��N{���
2Ut^�<ީ�˱��A>4Hi�k��NEk}O�m�бƙ6���k���9�?���@L\���gL��RCkX��ƶ�MMۚ��v5�}�a��c@��a��v���.�O�jw���';v�S�5�h�>��w�q��������SOL�?�����N��7eye��ڰdwv9���y���v횞����%Ț�B֎$&�}��«�,խ����D;0<Ȯi�;A��X��$W��H�<���2��Ǻ��ȵ��M+�?�z���W6|�D�k_]y=wkTm-�~��/|x��M�±����32֊�H(9~¡�v$:��}��	Y��D�j[��h��q��k���wn��y4����m�^�@érﶴ�����ӷ��ٓ����="_����7?�����G XrzQI`�j��j�V�c�	�V!�`!�"L�\/"Ñ�3"_�/�I��Q[s_���ky�t��˗�Y�|�J������]����	���K^���%?Y�Kk�A�p�S�Z��!�U�З�U�:泵g�6I��p�v~7�P�eጎk�����[?�=��M��)Y�_ߗu����d�G�u^}��Z�ѕ��:��I��gz�D[Q;��?>����ۅ�k�Bo�H_h�A��C�&O�j'����XT���(�z�Lr�\���m�)�މ�����"�V���3�.���i�g��n�wfκ�h�ֺ��}�?��P�kvD\�v��]-<`M�6���6�~+6��T��=��#�}��y�i��p|;m,V��o��Z�w�@�t���y�m�>|Ҋ%+Y�rъ�o���;cFͰ�WFn)>��ק�6EײAo��ޛo���Q�^߱á�ȝ���N��������5r��R�qA_.>��?f��FF� 
'��(��d ���{�2��AB��¬�,YS[�����=�5�d�6?���Vh����|&�v �%b>��Qq�̇����	rRc��j���JFYM�0�C�7O�ɷ�z�#���G��Kh����U��G�[�ذ+B��c�B0K2­��g�!�c#�l��c�9#9�yb��]�"�	?`�&O|���I���nZ���'���{����������m�����LF�K�X�#���\H� �v�X�y@�{��kʅ�N��o{�����׮_���׿�r�:��һ?��⻗��o�#���!H�ļ���J&��O\��xt�w+=�OvB,.��W��O7���F9�1�Y���"$����ҫ+���bmë�u]��e�k��W'��ݡ[�*��/O�d4a�q��7���4!�%� ǅ���&.�{`L\��8���I���Cp�s��Ǒ8:��?���cc��F�n�M[e�]�S��Ǘ%����E�x�\�;���,
�b�����~����8;�	6[���68$8�Sp����&k�	%pM�A��Ju�1���:Ym!LdL�7Ť�&u3B�e
<�ӡ/v���r+�ɎL�L��q�	�o�i���D3�{	��cj2>0�����ֽ�qh�̣���ޜ��K�Mڭ:uoƨ�a��/�}$,�X�~9�f�!=�\g)�2�ެ>	��䫚��!�OO�Y�6�b���<��]rZ�������g�t�>uj՛���G�Y�I�了�36�~�M_G�q����-��V+=i�l$�\k���c�k����ňS���-]�������g�3b�����������{�B�be:��yqݱ�"1mk�m9���NK���*N�TURH�I�����MH��v�	��� �r���,�1OZI�r��$�|\/�bX&��c��U�[��N��l8�Y-Vq��Y��<imMH����l��ѵ-�'XU��\#'mf��j1�c3��sF��xv���8ߙ���Wm�(�B;�����N�h�`mo�G��X��]�n
3G���� m���y�=ɜbI����7gY&�&��Y!�W
�Y�<�l6_�k^`)���c!<DC�!֞��z�Gba�h��
��l��,R����AЛ�T��a6v�T�ow�:��������9,��_�c�o�f�5�\]�ȳq#Զ�IS�r�$.���(o�s��-zZ�Z�T\lVh����yY��6g�K1kIv��������_1I�[�fʧ���t�I3Q�bmm���NR�[͐����.�L�Ki�EX_�Hk��s�;�Lo������e#X�~?}ܐ� q{	d 5qI>m}}��ؘ�����6�8��9���;||}�����$8Z�_K�锿��V�?�AL�ߤV�a�G/Wؠf������B́���^q�v0��9����O�o��@�����>���}P3�R��BR�5Q�sB�VO�X|����S4�?E���7��m�zZI��ȋYe.Y-$4. ��;�0r��q�r]�/�كW����^&�7Fn�qH��hi�|Y�j��&O(OXO:�Z;��P��!ё��Z�'�t�d%�Y���F��NɝL3�7ú�sM�i�OE���/���s0g4�P��׾�*�̀+Gƙ��N��W�I�kM��� �k=d�Hv�'�Tim1!HYl&�!~I�>Im$[��F��&�M���e �^d���/���S 3k�8�h�^P)�B�!r�|I��wY{�����l�K�U
���A�R�:!_�Q�P�{�6�I;��7����f���s���|�d)�<c�[�s%�|h�� �;�����y���;�o�cw�܁;p���w�܁;p���w�܁;p����"����'B�P���&�F<�6B�wF���6~IS��UW��T���%��u��k�u�D�t�},���/�vN�b��1k��N���3b�s׹W��UWI�m������w�LBm��ul{�]�ia��뾤��԰Ҳy�3*��r�;ccb�8g�s&VVT��eG:SJr���EE�tѫ�W�W>;/7ʚ�7+{|�3� �df^�3�<�YX�,��QT���--�.,����.�p�.-)M(-�|^yEai�36�� �x,��{痖`�JL_PYY68::��*J��s��K�g�E��UF�)��0��$7onTYAYtjaN^IE^�-�5J��V��眑WT:�{��W�e�6��N�r�Ƭ�~�e���u���,:+˳s���w�淤b���+/.���E�<�5�<��2/7ҙ_�1C{���Rgv�<gL��3*!pa�L̒�E�ʂ<�!�srJ���]t�, �"C��n�R%��A,י]QQ�S�������⼒��J�O~at�MP�����s������ܪ�<I&��Ψ�̓<4	+�U�
N�V�VU���B�D���J���@!N��8OJ-�[Q�5G��3���Y�;�w!Xu��bj�Ȗ	EW�U''�SPZ|� a����L�'�:+J#�U3f��T�C�EpI!PNiIn���b�՚�G�3Jg�I	/�4:AIi%�Pa�
��5y���YQ��f乵6�����,-�_�;�K��n+��r^Y^~6&�2�j��8{��_\�[�_(-����
�f��J�Չ��]������D�y�3K$3��T�A�C�s@�B���S�r&��r�eyhA�=��KE�XR4�Y���!Ry���WT*�2�m<K$~�g0��<��ڸC�ܞ�P�tC��`wt/XM�j� ��]Z��X��J�gvY�X���<����[� ��Y�]�y%����<<�Y�i��<����e+J��ʖ���v�����X��s�L��XR�?~�c5�
A,���F$9�Ǥe:3�$gN�OOr�d8Ǧ���������}h�sBJ�1�2����9�9&��6�9*%-1ҙ�56=)#�9&ݙ2zljJ�R҆��KLI�L���1��Ԕ�)� �9Fu�JI��F'������Ԕ̉����4A3D�c��3S��K�Ow��>vLFh$�lZJZr:fI�!@hؘ��S��ȌĠL4F:3���Fǧ������N�%
\��3i��1">5ՙ������?Z���6f��Ѹ���̔1i΄$����d�Q��Ƨ��t&Ə����4����Ib�𤴤���Hg�ؤa)�=��'˔=�{h"U�;lLZFҽ�Ѐ~�)`�Ir
��$gR�4�+�d�I�ldeBJFR�3>=%C���>�
{b��q�)����W�H����%F�LL�O���-}�]Iss��*�o��e(5�g��Z#����`�m�
�ʒ;���ؒ#��W�x7v##����C���T�9�r�c,.u�{�E��{!^faXE#���gC,+/Đ9兕&��*���wo���b�����U�a�*��W4/
}��~&9),AV�]�/�r�'�V:gJ��Z��J�!�.#�H9)$3I�$Nҍ��ƒ@�f���$�O%�J��#٤�D�5�����	�"���7Ҫ�wy��a�l�\���D�f��xR�9�*3eO'ꂾTJ���g����K1o�|֒N��"(�F���Rr?���+0�TҌ}Ȁf�=�=c��Η��D�n酄��o����\w����~���˟�c˥tQ���1�dx�%ZJ"����2�,C[��6O�G������c�[m"�U�/�v˃�J1[wi��5z��_���=g����>f�_y�������:A�B���y��j����h+��/B���^������,�-�L9K���\I'_>�k�Ͱ��{���R�a�_�^��'h*�.�^aȒ�ִ�f����Ȗ?h#<��M�CA�6x/j���Z�^^*-�-ׂS�`N��b�B��́WK*��G?��+b?���c�":�+�?36�D���b�*�g7�R�J�k3�R>����3D��R8��T�̑>P #D�[3Ų�["��f^ip[%u�eQ/���غi�V`t�O��(g��RNI�X�B�V�[���h�ඬѣ+[x]�Ds�>���Ր/#l�[�<�s%sDʫ��,�ȑ�>�~\䎒�ȹs%ǅnN�ՙ����224��;5i��H v�J�j�h�׳V�n��9���nK�h��_3�aD�쟱g�ܑ�n��k޿am�g��7_FA;���~n��ɼF����+�k����g��
��z����<�����W�d�q�r%��^%^ژ)�K���3ybh���w=s��O�/���r�yX����8�yN���R/��1�m�"9��g�z�;�I������T4z�gݴ�E���.���H�r����싡�r�!�{v�P/o3�Nj�}f�\��^�V�׃����69Y�{��� �.�-#k^�o�<���)���)�n�G�����.���U�,�[_�?���6���f+d����M�γ�DQԘ���G4�X&=�~��n��b��m��������R�p��J���ߨ�$I�3���N�3w�d��t�L�d�S~��h=E~ey��K�|"����8uAq'i4ҁ�h���^܍B�4�c���U�3$U�u������T\�����&�p/�É�F���0*S�1N�bp����Y�s�"g�p6w�?��4^�d��5QΟ,�i�|&�9��:��a�(Uމ�q��E���x)��m��!�Y�$�%���g�({���ϔ\��2�=#��B�D9^�:J���q[Yԛ�D�ui�!�?�q�)*�)��DK��M<�{�z|g��0�я�I�����3�E���ƞ�^V&�%�&8O�3�K�d�V��ֹ�wxf.�K��J��3��$�Oil1�1E�:̭[�����O�ziw��QX�^̚���x���R+D��$�a�x7楳&맹�;���c��ݪ�	r-&�^����ZH��w���q^��8��i䬹~=��������g��L�����0�Q�L׈]I��r�y���D�k�s{g�MY�w�I�b�w&`D��oq�~M�F|6���3�ww���sJ6r���ד}��8yg��2O7r��Ƭ��?J3�9�iӞn��e��^��א��=�%-#�̖ق���6�����	�L���,sd�ҝ����}E�������_��G�_���w1�T�R�"��r�-'��Y�N���[X������e*t0Ӌ�\�ō��ĜV������������#f"~A��_�g���g+e+�VԶ�m�?��B}'�/�w�gP��A�w�9����������av���˨��^A�,;�����*��++�7Q?��G�-�m��Q>E�3�g��_�`������?O���'\*��M����'7�����I"�˳g���y�E䞙�y���E٥N2�(���]Ej�%�2¨1�!+��	Rah��Z֙�;��Ĝ�1�I���8U��cR��d]��O�f��X�4RR�G��)q��}��/��.���+�E��V��1I)�^�Rb�mH0���B&~H�Ң��1G��:4����J���ƽ�IC�u8l��w]����rF:�a\;b&���.�@YY�e1ZyX�%r$�c��"�Ơ��cX�)T`�S�k:�Re9�\Y�,V�I��&�~�=zݧ�j�3&�d�IP2� �Ҏ���gs��?���/�OK��������J��z���,:J�M�2]��bo�:��څs�(�>�,��ZJ(��M'L%���V�D?�_�:�-�Au�0+s�6�#e�X���8��RY:�bSY.����l��-��|�m���a��^v�ղc�4{��g����+���nr�5n�<��.�������G�4��'��<��r>�?���z��o�;�3|?���e~��������k~�_��
S̊���W�J���*�{�De�2V�LQf(J�R�̇�V��ǔ-ʓ�.e��_9�UN*g�7��%�S�K�N�V��誢ZU��F����(��:X�S��T5]�R����,�L��.P��+�Gԍ�6�Fݭ�U���1����z^}W�P�\�J�F���Ԉ�iv-@҂�.Z-F���Z���MҦk�Z�V�����Vk�M�vm����O;��Nh/k紷���������U�Vob&���hjor�"L��X�@�=�D�H�X�x��:KZ<�����@�]���c���JW����s·�ix��Z q�����u�B*p������!�SGԥ��2�"�\<]/���Ԧ˖!�D�nz��˕�z�����T]�<��M�x?eq�A��^|��_	�^�+{���S16K��O��̿���C?�X�OwM���9+lx8Y�	��r�'q�l�W�,�2X��2]⥒r�ē]O Orm�uђ"�ْ)�ѳ�ģd�}�[�nt�_�O�L?u^)��>C�J����^]D�,�3e����KD�,����O��Vj��_ �se��M����1*�zY��&�[��m�s=��ʺC�Ta�E�b��ShL��?���8ȵX�������F]/ �(q�^-98Rh�!�z��U��CR�GH�#dK���4�o�f�v�zQ�v*��߬}��F]�o�ӣb�T7��X��pT�Ah8KwH�aF*�D�����A������t���ӫ�"0�*��^����zAc�C9j~�{��S��?յ�E�c������u�����
�Y�%b��N���

F;���K�{%Wb���OZ��-����A�H�{u�&�ZK;v�=��l8#֬���B���}�R<�/z2G���i�`��-�(�Q�?��+���1JG���hfĜD���l�+�L������&�
#>�e���2ݬ<MB�]��>�P{8)�w��$���w�9��02מl�C���"��'ԧ+�§�Owrŧ�O$�����ݹ�?��lׄ�7���h�ljע�	���<E���t�E�Oԏ���)�e�li�e,��ʌm��LyHY��]����d�+������/1�$Ư8�'�3�[�[Z
�LL�"M�������}��O?�����*�N�cf��Y{�d,�Ų����F��l<��f�V�*�|��=̪�cl{g�=8�bG�I�C�`�%�)��ձo��s�[����y(�ƣx_>���d���y��s�,^�g�|)_���6^�w�� ����i�?������W�~��T��)v%@	R��.J%F�Q�J���LR�+�J�R�̅=��V�+����N�e�rP9��P^V�)o+�++������u�^e�Y�U���S�P#�Xu�z����TǪ��)��@-Q+���b�a�Z}Lݢ>��R����C�Q��zV}C��^R?U�T��o���)�Ushm��Z��M���j��8-YK�ҵ,m�����ʴ��m��R{Dۨm�j���^�V��Nk�i�w��ϵ��o�k�M1i&�+mQD<�5�~^ub��Sj��5���z����pQ���EdG�:-���PE栈Qt�jl
����*��8ʴ����+uR�]�\�&v���NJ&p�*�ڮ�@�U9_���܊�7i�
ʬ����W"��ʎ*�.h������M|�\�[�E^�,�/�\�8�3��d�K� �t��
yY�ē�V���@QW~��<'(˖L�S��E�x�*N��	L׫B���5�U-N���)maV.7�ϐ�o���a��JN�d��Ļ%~��M�o"��jY��njg��h�C������ wVa�U�J.��$�&�I|S���,SY���V��~�G od�e����K���Eޒe;E�:VԅG�Ŋ�G:r�!�����|�]��?V
��u;?+}o��RY�"(�(�"��iYs�)W%e�'8�\��KO<_�N+��O>F?T�/(�1��(�%�I?Y����X��2R�gW�JN��f�I(���D6r���c��?PY)�D�opq���?F�;~Fz5�A�"����ή���� =˷�<���&h��8�t+�\P*E�"�FNhʕ���_����/�W�V�Y�� }HR?#(��j����i1R^��.�d����-�"��^UH]�v�Dz��\��o��!��E����O�A�'Z�Z�����Y�!V��+�X��\Xs.Qb�ę� zYh����
2"ī�h�Zh�����?'��7\d�˸���xw�ԋQt7L��oi���<EP�4�X��{��澨_^DW("S�s�0�I�a� ���S�S$'�I��t��L��g
d>Sd��O���d~�L&�|�����2��D�3�����-]�Xc��Nm,��.��a����F�4��&��,��r6�=�b��z��mg;�3l;(�gd/�s�m�>��]f_���:����?}y oϝ<�G�X>����H>���S�^�Kx%���y5�o�O�]|����$?����%�)����o��+�bUJ���tS����`%NIVR�t%K���*��2e6��TY�<�lT�)5�ne�r@�U�)��ה�ʻʇ���W�7�5�JTM��j��vQ{�1ju����P��Lu�:]�W��ru������Z]�nR��;�g�}�A��zB}Y=�����~�^V�V����z�if�W��kN-B��b���=Z�6R��צh3��D���k����j�1m����Kۣ��iG���Y��vI�T�R�Ӿ�nh�I1YMSSGS���)���4�gJ6���MY���\�,S�i6������GLM�L5�ݦ���Z�1�i�k��wM�>7}e��t�t�L̚�n0���]�=�1���!��s��@I�ʦ�(0�+��e}���/8��s����=֨w�}.7��=���f����1f|٫�W}�7���}����(dݻO{9���k�3�*�x3FyK�����m�O��o���7������/c�Vo�?;��V�C>�V���ݼ�����z���t��{I�k�ۚ��'��}ޤ����I��{ݫ`���ī�j������/���z��Wӭ+���F�0֣��xk��[¯���_�0ޫň��ҟo��zn��w��c���_��(dɹ�n҉2K���طY<���!�ޞ#�H��3�[�!�w���Y�#��R���%��2�l#O���Ԓ	�09I��ir�����ߐ��_H9��|�1%�Ęo�w�qr��@6����l%.����B[�]�mK���i��a�yA��hz?y����4�k�{�b�JmO۞�����Y�m�m��b��� Uml�����*��5e�5~Ҷ@H�v0aAc�5��k>�0�0�JL����Ŧ�Mզ�L[LO�v��������N�Κ�0]0]2}j��Tg��tä����0�1w4������}̓�q�ds�9ݜe�j�5�2��g����Wb~e�y��Ƽۼ�|�\k>f>m~�|����C����ߘ��oZ�E��-� K�����%���2Ē`aI�db��2%��e��A�C�Ր�X֣lBَ���}(Q[NX�/�s(�6��(��G-_[�Z��ZO�������(���V�5׊׊׊�
_�"õ����N��s[�s��J�b�b��Q�QCق�$�.�=(�Q��������(�P>E��Zg��(:!6�js ��ٰ�l�(�P�P�c��ġ$����mY���\�g���`w��OlK���>���߻�=�ٳ�	��S��)db�i��4I����Ƙ*���1�#ƈ1F��ҌC�0H�Pd�0�)�)�H�B�=����{��t2��/g�{w�9���{N��\F��kHz��i�&��Hېp�w�{��$�!���	��|F>��c�� _� �Hɐ*�C:�Ax�Q��(,�!M�#�� P�@�P�P	a)��UP�Pw������T��?8 ����ӈ�"�� u���ԝ�*����)�v��/L�PPs�x7aJ�2^�7G=%	���RPs�:��S)�9��~G�)k�:�AiTPg
�LiEډ�zSPo
�MA�)�7��]A�)�zԝ��SqTVQ{*jOEݩ�;u���Tԝ:L��Q'�9�T5_-Vg���
�u��\]��Qk���u��Yݦ~��R����ԣ�	��zF=�^Ҙ�M�Ԓ�T-]��2���(m�6Q���j��T+�*���Rm��J���i��F�I۪m�vhj{��a�vR;���.h�uIﮫ����iz_�=C�g���x}�>E���Yz��@�����j}��V���F�Yo�[���n}�~P?����v��~Q�b��DC7\�����g4Ì��c��cL5�bc�1Ϩ0�1�ˍ����Xol06��m��.c��q�8j�0Ng���%���L0M3�L5��� 3�n�2Ǚ��f�Y`�0K�r��\h.5W���s�Yon4�̭�vs�����<`6��'���Y�yْ��j�V��f���2��V��m��&YS�<�Кe�Y�*k��̪�V[k�:��j������i��Y�#�q��j��Y�+v�N�u۵{�}�~�@{�=�i��'0f� ME�GB��{m�^��F��{mUm�_��F��{m�^��F��{m�^{����k���G�p�g�B:��^l�;h�z��^�N���;�AN�3��s&:��\����:�N���Y�pV95�:����49[����Cg�s�9�sN:�����+��]յ��nR_�7��f���xw�;��s�Yn����r���jw��֭s�F��mq[ݝ�nw�{�=�w��v��{ѽ�NJLғܤ^I}��y�~�+ �B�[e��CU���s�:oUA�6��Xu:smg����#�S�����:��+�܈�%�� ~E��㭷�|����^��3�}��=�A�^� ?V[���p�]m��.�Q��ߙү�NK�r+���g]|��r[1K���K���Ϟ;Sf�҈Ϯ:�~N�z^��wu�O;�/�ƃ��yk�=盾x��T��W��Y�o~���>�KS~�_�g�#�m�uP������a�>G�A�܎���N�Z��o�ǚYb�����Bᛑ��L��)V[>�Bu����
I���������:3�ƚ���	��:�s��}=�=���왮m'~{�}��ʿ�fb�c�}��b��l[Mϧ�p�����T������F|�Ө�kur	S�;/�:�:�~��7���
��%�/Q�2�e�V#ğKr�?���Mu��d(�Jx��+I���u��-�[�[��ؽ��5�֧�Lo䌵B#\D�( �f�v>�5?�+�Ne��@���:�˭c�?�{��ue��Nr���F��|��4�i��"�B�Sb�9��������*�ʊ ��� ?F[��!�$�%�ѳ"�Oz6:��8�Y��	�!�Cx4�ф�	�.'\Nx�UҺ[��q+�V�#� <��4�%�K���㱄��I�g�����yў��i�)����b�C�?��L�ӛNu�. \���x�{~WB�$��������皀��.!|չ���&��i�g4׳����h��>�O���޲��f�l{����f��n6��agY%}��]�O���~�I�m��,�������&Y|��H��0)K��li�I��KCsCO�9��C+yE���^z-T�WF�"I|U�G�n�Bdqd1o�l�l�o$�M�7$T'T�7�Ox�oLX�����P�P�7�n�;�[r#o�ߕ�y3�l�݂����E���x�	���(_ˤL���RK��>��u7ed�GQ���E:�tI��B:�t��҄D� �H�H�H8���t>	�|8�(��D��D$ѓ+⚐pN�4�]|���H"ƩID�׋X �&���i�q��v�8�Zǰ��H��β����ҳ�����޲�,�Ž"��C[�ڊ��o��|K�H���OXOJD�b��2V�V�ձ�ȚYkE?������;��X;��Ev��y"׹�{�>���a|$�'�>���b>������/�+�^���|������E\hl,���煮�����
��c�oKx����e\2ʵ�GH&�Ǵ���4	I�Y�!"�S�G�W��I���h�Ռ_�LD�aOu\z=��c�P��W܌�����eѼ�s8���>3(�s�}R�g�}V��9od~F�y��)����4�gjz���u�0��1L~���i,g�c����,)/4��Bs)/4��BgP^h.�Π��\��%Y!��z�X4W���^H,�h���,��h�<�]\Z2���QR6�M*)+Y�� c�+�[T�w.�Ys����rQs�@��ѧG{�і#T&\�����)�_f�L���Al(��EsMgE%M���]�t��S�Q��tlGyx�J���|W�:)�WI�TtK���,R����:�jO��Lb�#��@d/��8���$����䷥�b�;i��Ƕ$�#�#ʰ��\�i�$Oȹ#*;t��!�����uR\�$���F�� ����ax�߁���0��L(�'`<	?���YX?���/�x	~��k��o�;�������#��(`@8��|���u�{���\�+���r�2@���Mfw�Xx�����Psa><?��s�S�9</�/�ex^�7�.xW�B�T����3�_ Ch`�W�'�o��⹆��8������b���A��X`Z�
��b?ֳ���"�&ڏ10r`
�B>B�CT�BX�`���P�P���B�|I>'�ɧ��H�n��)_�H{�_���
�A�A;�&�C�~E��2�z�V:ك�l؊g��X��f,�~�}:��μGgnHI!��,����O��
�z�Z�ا���J8���ʽ��bEl���5��{���O;��ޱ��?J�Ha
endstream
endobj
22 0 obj
<<
/Filter /FlateDecode
/Length 445
>>
stream
H�\��j�0�_e.������M�E�e�} Ǟ��F6�s��_YGt�q,}:g�L��o�~��zcw��N��_�[蘎|<	I���Y����NTE�p��|���H�5U���uwzx��#���-�����!��m����~����z>ŋ^��W{a������0�#��ğ��$�9���uj;�?3���4��ŧ!���F;���6��YY��6P��'�j�@n��p���� 4 ?@X( �A� �P � ��
�@j�S#� W��6eC ��
���έ���e��)��m��-�ֻ�hS�eY4�j|4��֊������j����e�FN�C{l.�6��=vU���h¾��-��p�����R`�r`�tY����`��0�� Dr�4����2�����B����;M�2[������i���W� �3�
endstream
endobj
27 0 obj
<<
/Filter /FlateDecode
/Length 14941
/Length1 35396
/Type /Stream
>>
stream
x��}xTյ��g�s&�B!�W	B��~���$$�2�LH �ę�����R�R�)E���H�q��Z��Ek���T��Zj)�3��^��d���~�~�e{�}�c��^{��3�3ƺ ��5mZ���3g�`�A(�==/�wbEc�ٸo�^R\�����)��z������N�y��[] ��˺;��-��h?����8���g�h��U+�\�
�؀�hssu���kF�_�X_�X�42�Վ½��nu��}�[�X�v�xݞ(�����S�����/���~@M}Ӫ{�������W�>���Y�2������U�qG�*�߀�w���'N���p[��4׳+1~��o�{��d$�;�Β����l��n�՝'����b��ƳC΄�����^�}T9�Z��~�z�h�v��<���(E~TYb�a�ĺ �eK
�!�K4�ה��Ƙ6R�n�����V����-tUQԏYZ�u�ϯAH�"+���0s�z����9���K/���������c����c��c~�V�\���ϰkص�)`kY5��nb����ǟ�VA��LG��l+���e�Y3��Y=�'�<��-b��nA��l�a{A� �*���7�*ւ��� �D�M��/E�uy�|l'+A��l"h�_�C_r�}���B�>>�T��UPn(�\ޗ�	�������]�3l�A��R�a��d���9HaA����A,��Zn���dA.�),��&bԫ�I��n����15�Zd�=�� �uH��,3�	� N�bD
���B������c��pʃd�`na����i!�&��A��%�����{�-�0�vAC�P�,�f�����&9ײ:��4X�A�ѕ,���L\����������X7�G�gY��؏Y�V��6�c�`��/)���_�%mXZ?֐���J{����#��gϚ��E���K��2��QB�zr-��%iX�U�.I�����@�;�<G��&]��z��4��P�l6+gt������&Ϯc��F�'X�6#U���zB��a	��b����(I�P�r��1S&RI���i�N@�L�<x��BOu�$�aG[ #!Eo����6��B��<���< n�s�y��?x����g�/�J4*O�~/@�e����������gr�^]B�Z�]�7�_�����P�X��A7�}��FY�K�����E ����k>�O�Kx�2��O���M�ݢĀ֫�3�K���|`s
�Cϡ|&{���;�=�x�3��%t�U�1W�C��oh�!��y���|,8׌��c�����؏����3]	k�B��a!�`Y? �XV��M�l%p�� Z�W�^+�|r%�3;��l�U���Y-K1��m2�I���p�W�aXͣ�������5���Ün�W�����c+Y=����,%��7��>R�Ah�	���f�6���mň�Y��ˊ 	h}�+�]�ǟ�h�~Dc���G�'�v�V�a�nvzO@ﾴ���4r�%��^{G�o�%@g"{�ƒrF�a��k'��cIߐ
�$O[io�ݏ���yI�N�I�J��;�M�|�ވ}'DW���H? ���B	Ԉ)�Z��"�I���r����m��2�-b�e���,�Y(��Y�Am�aƗ��G�^_��m<�m@����䰥�R����r�f@��X�{1�R�;p݁���H����sЧ�f��Y��� ��f���d��Y!�oA��z�Q�'����I�I����g����-��06	;�Aخ�8������3�DI0��u���F5|�B��ˏ�-�WX�VИ-r��}��?�e�ߌ�:�S����{-Z����r �D�W�<hY���G��R���[A�{\4����S��/��l$�G���@���C�{�Q��λ��|j/*�`��V��d��Ue��Q?w%�x���A5f<�j�aGC�Yv�����'�x@����d�M�惠�t�p�*� Ȅ�M���l�(FJA�x>�Q�5sQӝU�	����+��NE���Y�ȯ@�H.��z�t8OaE�>����@�t��L�BkI����:����0V$ET��Pr��o�5kEQ��!��o)�����\���D�TD��h�b�x��x�W/�H�"��"�,=3���U�){dl"#��$ǖ�Td�":+�� ��j�ֺټ�,��'��}�\�����/����uiU����������[3ZUs�9VK�g/a������[����\snDt]\���g����l�������\;6S�+�����Z�]�*���%ʅ��e���"�w��Ϳb��o��FJ>��7��}����a��cG����2����	t�A@^�XT���8��������"7x#V���7�0y���EQ�2~k��`;���l���6��X�o����!�Y������ r7`<��������*vJi�;
(@�xy����t\S��{�e<Dw\��o��`�g�3�y;��$�Yd�=��`I(��J[
?^�6�6���,b��t�sΈ���c�>�3��G����f8m���S�\�DVQ�·�,�~��R�'�d�bM������ھ���r�ѕi-��6��lǃ��pR$�B_tmOU���v�����
:qx U6>Gq�hW��a�y/X���A{&N�m�m����=�i�\�zXhg����n�ca}kώ=.������r�yd�gʂP���W��`��A��o��y?�P	�Z�IId�dB��S��j��v����g�S�(����r�}�H�.��bN�J��}Ly�3=x��;/���j�+{ȫ�Vβ<?HNn��1X)��f�'A�Q�ߕ_�#X�O�_�O��,������gX����R���X��"�J���yYo���}B��U�#x���u_���AI�����Y�j���.J��o���i�.����/ �*c��e��7�Ih�(U���cC�˼�v��R��t�M�8k�FZ ?;�<�����x��h��-�e�k�{�����nD���>�h���%����Ex�d�,Em/���p;v�î�=��� �T!����h3�MչX_�P� ��T��F��6��2ps�6K�
��ɸ%�Љ��j��Ė���p�.2AiNyl |�,���b�g��L�w�" �y&hAD7���81u�^5RF�`ȶ���Ȗ��(�A'�+0�C��Ґ&�d+z��ڼ	�l�>:��]��Cھ�_O��!h9��*�@s(�������vt6 �$�Ob���Y�pj��D
j��J�(��K|�#��dGA׏h}KR��T��:�%�2�-��'�KM��b-\^@�ċ���јWy���~H�jƌ�I#��e�қ5�t�
��@�����S�_��E��J�wɀr>��`wJ.�qw[�̓�K謐�����ʣ�� ��"��q��rI�|E��t�8 ��3|��)���K�#h�vm�.������`K��V�}�|�RW�r�Ȅ������]���
�C�Y�ay�Ñ?��B� q7�.1q����<�����y��S�~o)�¼�.;�/��_����38�<K|�W�C�AH�~�H�_���`�DǾ���h��Q�)/>f�|�����������!y�+�u�σ�1c�}2�&����{�U��߃��'��Į�Sv(��'�>������}��$'���� r�@��� 3<=��)]P.W�\�/c�uq(��r6b	/Vj-F�a=���W� ZX5U��U��B���g_m��=�����I��$y�m��HW�IFUH^�iHK�$#�Z;�f�$��S)��v�	i.�
;-�;����`:E\�����������i멱������&׾N�_��,��2ˆJ	��:��H��>�p�*�2\q�����9��������pd%;�v	K*�^ڂ�Z�"5ꠚ���7U��1���u���<�j��<��U +�P���<����R�`�AWU�뎸;�O�#�;a(;���n:j�'�O<)?'~qN~l�v�I��tq(K<�"�{���Ё��C�Ł�bW�)�������y'�����^S�}Z�������uꞟ�i{�=�����nS�4K��&��9]���	��Tw�$G�9]�$G��q��c��q��n�{ωm�ďL����a�hI�7�S|��M���mZ+�+A�;Qܵ1N�+Al�wV'kwf�;q��'��M���چ'ņu�m��j�-�e����[n���C��Y��"n4�z�[�%���U[�7t׷��q]����k�`M�X�$V�`�G�4�
S4:i�N�M��7�5����k�/I4�?�5���n�V���_��զju�E]��|�X��eO���`��A��X��R���H���'<��2E�)�k�S\���L�����0K,�E[�(*�|�E�o�yYb�)�˜Zy�(s��9�Zi��S��I%q��E�=ZQ������e��]��-����qNL?'���y]���"����$rb�YbJ��<)V�l�I�ڤX1�)&��Mh��9�����u�8�������+ƀ�1Ib��$m�,1jd�6*I�LY#��,���Ib����Dmx��$2Q��,�f�kC���G���h5cHg-#^dQ��ՆtC��q7X��Ǌ�G����j�,1��8K�H���T\Rg�P̀$�?A��N�R�D?�(���B�k���+A��S$�l�>h�'K�N�zv�z�"�F�ڳG�ֳ��i��#���#^��<�W�D�Y"�[D��"a��ʓ���D�,��şq����c+��kE,�b+D'��,gg�H��"�QC��,�,	��a��0ZյhM���}Hբ�v�����"��I����O���G�疻����6��Ӈ����~;�]ׂӼ�-b׊?�f R�(�H5x�٭��j��F"��D��$k+C�TC��'p���/����e�򒲉ak��MA4v �����BLu����9��s�D���)���c�xV)^��z-v�_q�ws�T��ɞc'�������~S��]�UlD}�#z��?$�sl���w�Dl�3�Q�Z٦<�.!�=N+��k�m섺��c��	�&�q��va/��j!;�^�mn $�'FkwY ���ڛ�d���%��$�pJc8���إ��a����`8\㤡��E��v#.t��نz��Gy�V��lر�F��㧎��5�_|j��~5*;����lqĞ�ү������'>�,N�{����Qq�_<�"h���b�p��Ay��Z�T�Ȅ�jc굠a��㢣�yk1z����zw�;������G�lg�CA+�ǩ�t2���g�G)Bq`%�p�G+
O�N��~�S��vA�#��9_�]�9�st/����LV���"�6e��㡘_:~��]<]cq�'���u��I��.z3���'������+j�����p��=�ųƔW<��{԰nܸ]������ǋ�"��<�䑇y���/;M~����uk@���r�+�>�k���Ώ��Ae؋���[���k_3�p���u��?TSյ8�gf��q'[�X#:�i�����]�{vM4�X}tOh-KN��3�Μ�;���ᩱ����Ǳ~Y���3y��[B�Ȭ1c�ԙ�*�V�]�����˲T�i۶Ms��?d�x7>~p�yf���{�?A����DXh��c�����Z��Y�P叽�7��*KT����}h
��F�a�NJn⻌�?�&F��%>��ȬDN����Dw>�|w��O��on2w�]}uC��W׉g������x�͇/6;�:rd��k�Z�Ք��Sav�[��;Y�M��k�j���$RS�n��ȌM앨��w����u*��q������W�W:��J�Wzi�������K�Ru���P����0?6Ǔ��O޵5�o�����J�ѻ�9v�`���x>���yf��7N���6�����
u������A={}����>]����,j��>ps���IO����.z�+=L�tw��Ik�C�Ւ���qz�������d�������ŋ��f�b?O�����C���_y݊!wW?��G���Jn�c�~���c��Ϳ}ޫ7�|��"��9�㸅���m*�.}=�f����nFL�&�YW6�T���q���t���IǤ1���/�
3��c��������+��<���T����O�Pv��g���gl�K�(�I4Em��rF��
���?^� �1��'b9�����)E�����^;��KN|�˛N�m�P	���~��;��U���j:��͟��%S$�Id͖�ĝ�Cj��r�8�X���ԮZU�lժ�ͼ�g�y��ӟ����������;���s�_��Ɍc�a�d���	�	":�%���ۍ�1����$;%��>~,�ZD���nr5u��弪7_?{�iI]�?��!���%�dd�LI�kh=�.9���Oo��~�;cd?˞��Pb�}���GLr����5ƙ�W���LX�T��oԚ��������}{9ؔ^��c�	)��a�?u�p|�끗���W��-�����lq�s�JzTztzL�3�H���uX°n�����'��Mw�7``��<��*ɼ[��?lژ�a���Qc��ޜ�**=o9�w��Ó�����^�t٬��������M�d�F�W�%�~������l�I��MJ钶kîC}��c���ue#���XD��X<�l�6�ĸ.�	Ҡa�Y������m��ms`q4Y����\_0��W�1?@���|�D��Y9'�{GQO�)�c�W�0��f��(�T��v9�\�&�f�3.vI6Bs���8�d��c��Eىv�
]�|�B��)1LB5�l���.У�{Es��^\]on7hn���.�z'^�XZz7�9�P��1c-m�v�htO���J�KS������"�{�1f���{M�יGͿ[v�$?��������k||R��7?�8���u�O	C����<�/���g�A�Ew</A(b�xA��&\��p.�e���2\��p.�e���2\��p.�e��'��2\�K=�I���e{5��[��pg����V^�n�r5"�1�5�y�ue��|�g߷�Nև�󝢿�޶�l����Ѹ;���s�r��y�E9g�y���Ո�ƒ�ev^gi��(�����w�	�G�|��iF/;�j��N�5���.�ir�Jwe>�U�ڕ[�h�{������LWN]��T�
�J���ד��]��쪪q7,�\n��U��jl����ry|��چP�2wC�5���s���<��@�����9r��@��ꡲ��S�k�pM`����q°a��h����U�j��7���4le���a���ƚ�a��Uކ�w��<I����^W��η2=��$Ȍ�i���.�rXo1C/�����5��0r-Xt5��o�ۿ���H%&��믯�vѺ���b��~wC�ד��Cxt���^����r7�v5b>��W��k�b�*0-[6�x�pWU���\6h��:KӮA)���t�܁���֍����zoC��I�S][�����Wݴ:OI'N��F���\�%2�ZV[���%�u��,U�5{$'+k�j|�M`���H��[��� �Kq2\�^���7P�1F�s���
x1h]Vm�;-��F��&[u4��_���4T7�0��:z|��/�h�\�j�%���`�R�*_��V��S�*w�o��$���A��	��J�4�Y�U�
Ը!T���؀�����k�]�]�>���b��V7z��(�b�}m�{��_���V�JCs�5���Q��C�[�����_�un?��j�6K�V7�d'i��*	�!~G�,�c)�]A��_��6�`��n�����C$�W����L@*S�Mh�xaw^K��>�'�J	��9v�"�n
��c{'���$�6c�+|�aƼ���j\��F,1we�WVX�r���q7�j�P�6���k�p��.��+��_I�$�������i��D�]u҃`��6�����B0�E�������n(8-�譫�L��wM+.*w�O+��S��*(s���+���s���>%�5��|F��rZ���/pOs�-p�*(��p�W��旕��K]�K
�QVP4�pn^A�tW.���
f��hy1u�I�Ib��K���mNnAaA��״��"Is��JrJ���-�)u��--).��<�-*(�V�Q�g�C�Z\���`���t*Ga���4'/vN��a1D.uQ�Lp	��y�sٌ��BWnAyYyi~�l�VjgzQ�l���Ey9��E��|���[�o�Q����p���Ι�_�6�lf�Ӧ�az~Q~iNa���$j��@���S˩%tM�S������Eڅ����ȧ! @�M%�H�"�+����Y�_P����)-(�,L+-�r>�C�8���Wd�+�H�]hh%{�����`�dザ���UU��&i����#�R�f��ZN &<��*�,�+�v�õ-.�%g��W�X7v#��zVx�ҕ`}��3YY���m��g�{wC�p+�Kw��l�_P���_�.+��Mp&.w3J��k��ooU%��t���4b��]�[���~��'����m�I}UMB>�ɵ��{ 8b�LW��|�W3?�eKY�gĪX:�Yl8`$r�h�b�h��H~楗e���5�}&r9�G�.V��;/�^�'����ay�-�y�-���*K��yI�*�����:�U��~��B�u�SFT$��hՀ$y���-$���,�1��mG!�?�{h�w�q��ޒ��ք��	�N�?S���W�}&��p��/�������&�^	��##�d�U�m�F���^��˦E��Sh�.�Y�?��s�?�\��r��k� �^�u��-������B{��?��WA��?aîo���֢���4�����(����)Y	ѫ'jm�kѮ�:�-�R����Ct���͚a��2�/q�@���a���&{�k�*,Y�lM�h6�W����Bm�!
���{];����a%)4snZ� ����m�g�`����4QMH?��G̖
��6����&����m:�%��>��L|�q�!	����KC��64�7��a��*p�LT,��$�!�dk���"%
����J��f�aF���|=�gh���o �3�A������K����,ڵ�V�����i��1l�M��M������4Bh5T��m�%�F��!,�Ƞk3�����m"��������=�q���Z��v/��=y��9��Em��4П�[�!Юmh�4^�D�s��n{�*�~;dk�6,O��|�hGr�s_OW�`�e���o5yI;���.�W�du��zZ}���CM��d{=����M/�j��H��_rK_͠�~!�<ĩ���m,�=�]8)�C�d=���訟�����<�,�Mst1.�I��:��b<f��^G�j/��������Ja��������w�v3����P����)a�;���C�nJ��Yk���>SI���k��B3���ј�ɚ�F�nX���<�7�#r�-�/�bj�ӻ��y��E}��X�]̇��f;���W�%㕔vs���ـ-�lIB�.��dQ�A�v��ɢ�/�g���h�c���᱾Y�J{�4��buXS��r�bV�;9N1���|ē�T'_t��C������P��O��8yI��^��i�K�P"i��^��B�"В}�Y��O/T�-K��l��o��=�k���^�3�Z��W9��O�bqZ��Q�sU@#�8���RПa��vѓ�g��d�(��4��ґ�,iNG�t'K��Z�ve����ⶈd��zK�|���	�����`l�B�<����#��-3HB)O���΢R��b{�e��J��K���:?lR~��N�_��r������t�0;lGsI��C1��KuR�R��ᖥ�2��%�Mr�G#�F�.*I�Z�ٹ�u�F�N�哦
�u������H֩�n-���[6Q�ݩ$���95߶��]{)�"�o��O��Y��ٳ;5<��deje>��|j�Cs]��4Z��m��FXXh���Y欽~C�(����Vh��3�G�ThsX�Ʒӵ|W>��*:�X����w���-*��?3X����,/<���wh�Vj�gk�j;�D�p۹B�d+�o�~Cч廭�Qd��8݊���?|��d%ն���i��ZD��4�%Y�ݣ#-+�tS� G\D��ڡ:�i��FYI�&;2��5�me���b�Sշ�AH�oӿ�滑Yg�ZҰ�'3m�~:���Dj��.��ì�Y��6�u�C��Fp�g��^M�c����������LaQL	�7��2f��Ma��Pnc\٠��m�6��U~���Z����ۘP7�� ���*򯩯#���>�'�0���y�)�?76�0�x��FR���19f;�>ez޴�r����+����:6e�߻��Թ}.����� ��$M�����S�A�0^V�K"���#\�W�(UP6��F�"\Hxvq!p����lT٬2�����|��zN#�Y��~�l�1��{����~�9ɒ3�%��l �v�wU����}��0��盭��u�}�.��w��Ɠ�[�IO�7KNaI˕e���>ꭄ�S]��!�ƒ�����Ԑ�	�oI�7���*��u�MdC�.�/I����9���e��A�#�AΞ�(�2��LaG����}l�\L
��
�烗j#�\��.�.�>t�ݺ.\�܋�Q���ӈQ��bP��,���׫롣$綮�GK�ˎ����/��~�����芡tQ��de�2X��Q&)���H)W*K�j�N�+��땛�;��J��]٥�U(��'���_+/*�+o+RN*�*_(_)�"�D�H=�K���%Ɖ)"O�%b�X$*E�hMb�X'n��U���>qPO�g���eq\�#��S�KqV���ƨqj��[MQ���(u���NS�R�B�J����FuV��X�w����ԝ�u���zD=�S_�*K}W�@�D=��Q�i�/�����%k���pm�6I��fhEZ��P[�Uku�_[�]�ݬݡm�Z���.m�v@;�=�=��Z{Q{]{[��vR�T�B�J;�+z��'�=u���g�Y�8}�����K�y�"�R���&}��N�Uߨoѷ�;���>��~XJV^Y?�������ҿ���Cu�8���ގ� G�c�c�#�1�Q�(uT8�rx�����0�O� ��5�d���5d��LX�2)X\\ƓZa�����:ء6��]��ֿ�	�%f��5{}�����V\��� <-?�|���^��w���j# �����C�A��jk�p������)ѡ��Y��Z�����ߵ���d�d�W�)���w��Ef#p}��k��V���h���$���ǔ���(�[3e����'���(�T+�SQ.$|e�^���픗%��SI9a��(³�d���x���	f���y����7��+	7��;��Cֶ����u;���p�fs��>9zD�c�4����D���:�JFɱL�bXYG|>�� 	+?f!�^0�Cyy���H[v�Y��h.��]�W>Ŝ����~��9���D�\l#�-�i�'a|_p9��\*�p�9KzA�&k�gԫ_�jI��[�Kb�w�1�J'�&�xi���|A�N������W����+/�_k����VD|5QXL�GTr_�?��9$�߃���o�m����Tb�?#1Jn�s�s+?9�|DDy*��������������#g������.f��E���^�Qj�C����}�k�,�s:07�I��7X,k�V���b*�.5F+�kJ������?�6�I'HW?��Z���W�c���H�`�Kk���גg�$K��$Z/O��?#�P�by�����^ʮ�4��x�(4b�Q��r]Iq���Y
bLi�7Ҙ�H72X��dLb+���=W6N��������d߷#��/�l�et�cn��M��%U�sJ�G��P�����-���>���՛ԛ�[���͛Ƭ�%�_�4)�Y�Е��3OJ����A�1�[���n�L��A���q�MEŀ�3�S����W%J�U���KIS2�,e�2E�Sf*%�<e�R��(J��FY�ܪlT�([��ne�rP9�<�<�<���W�Q�W>RN)_*gS�"FĉD�[��A"S�D��&
E��W	�X&�
q��Qlw�{�6�S���#�8*��ī�-��@|"N�3��T]5�.j���P���1�$5W�����Bu�Z�֩~u,�f�u�ڢnWw�{��!�	�i��������ԓ���W�yMѢ�X-A멹�4-C���iS�<m�V���i�Z�֠5ik�uڭ�Fm��Uۡ���i���Sڳ�����q��}�#���vV3uU����D�����3�Q�=[���z�~��ї��
�:�F}�~�~��Mߩ�����G���1��U�-�]����~F?�`�a8�8�Ɏ����1�I�\�G��ܱб�Q�s���;nv����hq���%��(�#���y^�giW���<Q���5��T���6x��<�_�}���S�n�������(Y� ~Tw �*0_�Jϖ�?'��)��ZW`�.G����]C�uY���L�eD4X��ץ��o	e�r�4U�<������b�Pr�T�)=d�Vܠ<ׁ����z O�����!�$V�T�9׋T�/�O����o!�M�<_Ix�\�K_��h�P��
�p�&�;��|�5�]�ɓT�&[&i+���p�Q&j/�����Gig��i/�rȨ&VG-wi���4D��)��~��]�C�<�'���u���*$?�E���LZ叨u��#j�,We$�k�<\~L�M�2B.V���&�L��5i5_�R��U����!��j���3��TrFbG��Z]��-�(�S*�X�ߦ��=Ң�^%c����dM�L�fH;Q�j�RK���j]�ܡ?J6&)�$�,�R2��7��d��mJRT��VGJ
�����&��<��=��Z�m���z'� �r��Lk��v�ܑǨ7��G�QZ�Zw_b��(��.K�'օ�*!O���r����I+��qD�!�*�G�����a0�1�3u�w���Z���^/�/�����ʘDW��x�*�
�S��ٟ�:Fa't���]rrR�퓫�}��B�r�?�!6Vb$��	m:�@7K��c�5	�J~�MFs��4S<��W�Wڒ.�i��J
5����>w�����H������]�nϐ�vH�BZ�����P��M4���+���7H�{Tɧ���.!-����a�pN"u��A�d��͔�)yԇB�TI��ٗ��?�K�xX�g@���l���4
g���|�ED
N;�Z��P5�"�k(�j�j�q���������8�S������2�W��Q�G�q=3��cxO�_J�3�(>�g�i����
~��e�������~7��o�;���?���������/�N�[c��7��Q�c�!���65�\X{!��\���Db��G#�K#�m�Ί,�.�;�_��w��ޑ�E����%lIji�������.�7�G�:��=/EYԾ@^�O<S��p-��x�c��`�o��]��A�=��}h���}��Zg�-��K�ɛ���-�_�� O#�~$�^�(�7�hn�Nl�|q3�sy.�@��=���_c��G�#6���ɦ`���e�s��UpFfSq�8��>,_���M��ݬX|_�ü�>��-ultld��M�Ml�c���1qkp�u�e>�>������A�wt>��C��X��M�[l���l�|#;=]a�\��F���EH�H5L�ʣ��.k��!݊�ic��;�v#��D:��ҳH�#������4��Y�zX;Y8��L�o��<��Zk ߭�m����A�Ð�Y��2;��aﳏ�)�<g�3���|{<�����7�����(�K��ғ���5�E˿��w)��|�X�j�����=�R����~�!.b��yH3�]�<¦�mӜɿNFL�,�RmD�Bԗ>xqlq`�q�c�8���}^��Yc=k�F�+�Yc%=k��xj���Q���9��^�g��E�N�_)rN�)w������9������@V��
zYIO +�	d%=���'��'�<̑U~:]�x�8O]�R6������jj��L�YI�����#����e�~ٲ���Sr���5=[�ԉv�ߡ��E�gZ�f��Bz�)gߺ�c]�B��Z����Yk,e��O)��:ߢg��	eS�ȧ������FĩS�l#��3�3�B��(5����J�ڨ1�uF��7Vk���[�;���-F����a�2������9�Ώ��:�r�6b݈5�IF��4z�� c��"��^�@��T?��-�7>3>��
�h�0��r��Xd,1<F��d�2�3�7���f�c����i�6�������3�O���g�_�e�	3z.#q�¢�E���z�z�w	�ȊZ�(�Y]>��N���T~�i�1ݘm��+���*�g��Ƶ��M�mƝ�&����{��?5�79�v�����/�8?7����ltu�^F_#��/��Y2�X�� �L1fRS0�v��� �5�X�`<��<�Q�l�a�)��Ts�j��6*=�r�P��X��C�B���&��_��8���w���'�zE^�x6=κ���&{�
endstream
endobj
30 0 obj
<<
/Filter /FlateDecode
/Length 281
>>
stream
H�\��j� �_e����n�B`IYȡ4�$:�
��1��}�	[���ϙ��3��}i���>�z���:�0�4�3�J���)���n[<έT���\���p�f�`�N�Sz��w��VkpF��uǐ起o��������W~;�_��f����F�b{���Bu
���V��?h$ɆQ�z�󬎆_�ɋd�G��('z"�D"
��g"JV�%�
]r��{Y�WR=N�J��)YY�F�ǖ�����saT�{Ҍ�t���Zc�*�_ Dg�
endstream
endobj
31 0 obj
<<
/Filter /FlateDecode
/Length 1134
>>
stream
H��W=o9��WL��H}�{�)���8���9����ő�d-i�N��I�ף����#���<iܬ�s��B����	f�|�:=Ӂ�Ü�l���o��x����CpJ[:էѿ���>w��#��>���D���S�9X����ez�5:����՚��.��������%�M�����zRX���M��d�����4{`�v6���8���Mt��ʃV��|fo���㜟˷�>~�8,���D���p�h5�w�<4p �O@2`�YkDΪ3�2�ia�W�ȒS����*��k����R4�Ń�_��Y�#
*�Rσ_+�60^�X��E%��)^����E�|��f9� "���B��	���^�#a ���cA��7���4��i������4p��x7�P����ĂЩ��UFr�z������y�������� �Q�[f���"WeqD� �-��HӢ���ꢨm��L�m�ΐ�&	(�.Ë�eX]���RQj^���n`}�O�/O6[ ?�T_��:7�ͼm�#y��)����%P��Y�M��Q����������Q+6h
p���XT���4p��-��M3�wlSK�qĠ;T6��������}�X����P�B�����6IWl�zv�qz�ѫ����o)NGr�=�1��Ч�;��l������N�|xҢ�]��λ�r��+�g��>�D�A�I��qh��"6Y6�ߠ��,�K�E���$�iD�Zp�����g�-�(��u�M3d�ְ@,{;R�����g���V:]���dZ��.*����	@n^@��tN�\�G��MIsG2����,*��|'�9��y�s��Wj�Q�'�Oh�}�v��.M�B��Q�o	�k�[�D`�{`[���{��vʹ;0��gM�vu�%�O���Z�b����μ��0���5W%���c�6�X�C������n|`��/�vi��<�қ�K(�!-H��-�l���y^�LfI��rN�P=b�G��ZT���r�;� �@�>>�1���b2k>�I��\k)ők�U��iP��Y5ܮnA���&�ۖ�!7�}�:\�A</Ӌk`�R���m�Z��^T�R����n��i�Z)���0�/� �ړ
endstream
endobj
32 0 obj
<<
/Filter /FlateDecode
/Length 927
>>
stream
H��WMo1���3R�=IU�&�7���T�����xS���J;�C%q6�˛73ϷZ������p��'���5=n���`��4����M�����G���Q���4Y�W���2Ni�O������f�H�k�.Q(㕅S(�����8y�(��N��"��V~><M�$�}�hkTZ���e5:��p�p�p]ᚆ`�'ES�V�RP��Ve0*�	2Ў���!oT6�w"dƪ���V0"� �����U2�e�:��m[c�J��O����MT���"=���Ç�q#��q�wjQG���)�ց�B�	g���(�������I��a�f8�R:]@���*xO����_�ti}1���u�����҆�����d��_YJ��UJE��,�2v&���F�@I��)�&�ۨ���k:��H��F�&(��\$y%�?��.�w��u1�x%zE�zf?������*��Z\Z��D���P�Ep�U���Sh�S@���
����=-DJ�	��4/~.�W ��P'���+6��H�@���D�Q�xp�&�6(��ŷ� G�)긮�q��L��"�N�k���3�O��ٓU i%��α�&�%��U�þ)Ԝ;�IkՐor;z�u�Zy"����sr'[¢�Q\*oY�u;�_�������������Ň`�s
R�L��C�-�ř��t2�G�̈́�2̄l���pd�z<���h�}ujG�9���]��Y����-�g�N�^>C �RW�Jl���23�^ n&U�KVtC�b���	�tԁ��ޮ�Hs�̋+N2.i��VB�*���@*��в�ᡁ+�f�?0�T$jc0��m�Va����תd�����i8�5ɲ��xa[��6�:n=�U�N�A��V#HM��^9?����  z��
endstream
endobj
33 0 obj
<<
/Filter /FlateDecode
/Length 681
>>
stream
H��WK��0��W�\�A#�^P��Ko�JO����a��ɛ�-;��c�T�c��<��C8"���||��ͨ�mƯ�!�:��8��^,������1|>�q�Vǥ�a娵���<|~/���_����L������Ëe�pK����<��2&��E�l��&� L���卓��"8Z",>�H���u���ȿ�h�e6�
a%�Q�EQ]�UnƨF��_:ZM�)��9�)�KJ�l�U�c���������6AGT�fx�P������XB)9M�fA�VNB��ѵ:�Z�Sk>�	��3i�|�diX���^��挎FN�@#@&�?�^rU#*b�3�ۯ��1��Udf|*�S�P;5�ټD'0�%�s����cQ�Nh�.b���8Y�l���P�<�U�H�	��q�pw��)���e�Xi��^�!�7��&0�v��Mx���K?�*��[B�g����;\����B��d~�Qx�R6C��@�凊�Ϛd�����1/�2������%��@<,�n�<�z¥�`��9����$AW��	j��{&��x��B�zZ��&P���$���8ސ��J:-�j�]	1x�u�Haj��� �~��%�#��)dj�;[�l��p����p��K�y��)L�ƃw_���#��^��l<��� Ǣϋ
endstream
endobj
34 0 obj
<<
/Filter /FlateDecode
/Length 779
>>
stream
H��W�j1��W̹aɲ-C	$�z+��ThK���?���3iX�[R���xg��gYz2����E�>Y?-t`8=�'������1}&��w�|�h�H�ㄳ~~}��MO�t:&"��y��n����hӔ�@x>���{}�1�����{gJ�� ����SB�n����9=�m��px�����EDFV��Wא�W�`6��n�1@��9-4��w��P��{� ׌W�V�j ���:� �^� �C�� ։���%(^2��z��lb�y9��L�(��0y���<�!�K�i229�� �Є,x�}X!@cO8'�q�G������2�L[�ŘO�0�u�$ڴ~#�R8.���͙d�͟�3_,�9�Z�g$qU��eo4�2����ӂNӆ��3��ۡ2�����sh��Y�Pa.�h5������vw��;M�Ϋ4�x���tV6@�]=��zT0m�ȹ1���}��m�[�Q*�}���j��α\)�p-���z�N�M���K�h�2�ѯL�)+�<Ǡ9l�sZhV��k@N�G��+]C{?@6��o<�!�u ��c�-��U�M=n���0y���<�!�K�i22�T��&d����
Y x�9A�<Ҕ����e�����1��a$�	<���o^
���9�l���r�}i�����j�_����U=û��Ѭ
M~)�\��T��%r����A�����k��}i���3\�&Tn:����ᦫ2T0mV������M�����  v�ҽ
endstream
endobj
35 0 obj
<<
/Filter /FlateDecode
/Length 788
>>
stream
H��WKk�0��W�\Ƞ�^Pْz+��ThKI��?tF�ÖM�H2%`��Z��ӧO�������(7#y� ֏�?:�0X�Q3�?Y���{����5��0|���` �<�Փ�T������_6-�L����1�^���7�sQ����-�$Ӗ ���
�t7�W��Q�$W�8��v���E$&� r^C6..�l,�	\�S���s�hV���a��p#pɸq3����ŀ�Q�:� �^R�C�k։���	3�ɺ��[���,(&3c��4Lހ�&6�@��]H�1���R�8T!l�d���"� �Ox�!��ͅgꄗR>m�H$��ExV��oO�8!S�5f����3�j�䍷*#��~�|F1�����DUgHQ���4��{��i�M���m�������S]�1�w%����0'�s5y�;��w�ӝ�u����٣pӖ=��R�mf�OM٣�is���l����ݶ�u�e��m|u5�.j�Un^�ẬCL��R��f�N>�g��K�d4��h�L�I+�<� i��4ѬFk׀��\2���h*��y-;��_;�N��7�b��
�����:�7้�%PAȱ�>�Lݐ��!e��C����)�@��/�N�Qx�!�����3u�KIi�G"1�.³�~Cx"�	��1����ŘiWe �z�2�����g�*��m��hT����^+nke�ߢ�����T+0��w������]�Ӱ�Rk�<�^sG �۩��R����qn
��{�����  �ѣ
endstream
endobj
36 0 obj
<<
/Filter /FlateDecode
/Length 785
>>
stream
H��W�j1��W̹#˲-C	$�z+��ThKI��*y���3$���2;�Y���,?I0��89k\��ٲ� �\����O�W�<M`���0_=[1���q��~����䦿�#F��S4y����鿻lX���h�|z�>��>���N���Dl�vA�'�Yk�I�^ ~��������n��ⅷ��O_޿��^B4Ly�xs�� B�p��Ik��<e��x����{,��_�kI.W�pyD�袱�`<��3�D&�� 	���78_ c��dA/B�&��.0�z�\�L�� 0�N4
B���&\1�y.�gH�1��8T���ޗm��r4�@$�#��N�u�I�q�ѫ���^�H�����9JI�]rr�s��k�UрzH.����}T�����R�B�rrB�]m[�R�U0�*̳5�f<��w���Ne]jz���G�3{x�A��#te�
��uq��5z�w��֝��ۡ���J�z�V�	\Y��uUgmҡ���7Etҭ\\��m}�M���j���%̅� �S4i��$�t�Y�ޖ��45�˞a��v�6};��_��Df��Zvf%����n[c ���%����LÐ!dIY �؄,m�"�Zh���Iz`�J�*�ߗ�m����4�D$�C��v����p<#S�W3��-���nC3�/�^4*��O>CN�|f�Z�FU5����k��Mg��X�{�V�]�rs��pw�;��>�;�� ���٣vә=�&)�7��d���%rn�5x�?����  �c��
endstream
endobj
37 0 obj
<<
/Filter /FlateDecode
/Length 791
>>
stream
H��WMk�0��W�\� �F_Pٲ9�V�[驐����茜ld�$D�R�q4V����񛙻��&�Ί��G�G���Oz��Ϗ��??��f�������d�<�����-(�'u�~Nw�����_2�6��lxe
��~���2ק_���Fp6��6pgli%^���g�_����
�����|�l���o��o�DT�B�	����������9z�<G��f1^�V�9��7 ��+��I�|¤7ZXG�A�[��O?�:A�?=��B¸X����|/k�Qe�b[�S਋�5�h�]�%�!C�$e��|2���E`���	�@"�E���ӷy੶��QhG"�!�g��<��������f��\�jr����.��0�*��c�و�"2�gtp2�P�tz���D���4�����b[��XۭAF����5�����m��{{�Dȹ]��/
7�	C��m��+c0M��S'���Ǽ��vW�MRg�����Wm���M��:N�u��Q^]G��ɢ�|�l¶��:�T���/E5a*E��,Q���K4���&h
����u�@e�@��@ދ��4�u�~:�u$^b���`��\nj��-��)p���h��>� �Yi2TIRV��7!�L_�<���$=0�P$����y੶��QhG"�!�g�8�F�q8.����L4<�W5����&��Fe5�]&�a�U>�ǖ�U�(�p�Z�p�W+c4"����V.`^�%����vw��w�Nd�y�x��Q��������+{0M*�Sc��������
0 �F�
endstream
endobj
38 0 obj
<<
/Filter /FlateDecode
/Length 877
>>
stream
H��WM��0��W�\Xa˖?�,ta{�0��S�-e����JIv&V�����i2qL�<�OOv����kx��_b�"�?��Lge֌O���W�4�=��0|���a0iz�4�ց#&�'��1�������|��2�y
lw�Q��u�Nئ7�k5�,��A~c����.�1v���GZM���~�r�Gd&m>"B��7L�w?��|�G�><�y˳�E0Σ*�}��״F�zM|�I�#T��C�ft���l��7�6#IH�y�6F-CP$�Yq�u���W�-w�h�ۃ��mS�Y�%2��%/����i�����I�6�����)g�R��B��)���%�Ǣ���-2#��;��2٫��Ƞ�^Z�j����I5��Z����C��b��8�ǚ��OS9<�8�����5L��b����������۰!�k�CF�������[��m��2J��P�W��7�O	�v��W�m� N2�׼�_�$[GAC'�@�ͣ�v�f��HK��ݢ�|yUj��VT�;�b�RZ�3P�����',i+Z�gj��T�0�Gן���v�3�����²�喪6�ѢX�k�����${}���u��i�W��[�^��9����*Lc�(�a7�CS+��^�[���i�[͐�����i���PjgC�!��4��y��
jɭ�%>pm����|��z;*ց���z�D[��Rʠ�[�S�ŋx���4�$Y��S��"E���L�0�LX/�2Q�v���g�'K��$��藆�A��vB�\���E��<�D��V2��Su��r���٣�aI7�u�<�_���_�r`0b������DV'�/[0
q�R���c����up�? 4�ű
endstream
endobj
5 0 obj
<<
/Type /Page
/CropBox [0 0 612 792]
/MediaBox [0 0 612 792]
/Resources <<
/Font <<
/C0_0 6 0 R
/C2_0 15 0 R
/C2_1 23 0 R
>>
/ProcSet [/PDF /Text]
>>
/Contents [31 0 R 32 0 R 33 0 R 34 0 R 35 0 R 36 0 R 37 0 R 38 0 R]
/Parent 2 0 R
>>
endobj
2 0 obj
<<
/Type /Pages
/Kids [5 0 R]
/Count 1
>>
endobj
42 0 obj
<<
/Count 1
/First 39 0 R
/Last 39 0 R
>>
endobj
1 0 obj
<<
/Type /Catalog
/Pages 2 0 R
/StructTreeRoot 3 0 R
/Outlines 42 0 R
>>
endobj
41 0 obj
<<
/Producer (iLovePDF)
/ModDate (D:20220227153102Z)
>>
endobj
10 0 obj
<<
/Type /ObjStm
/N 19
/First 142
/Filter /FlateDecode
/Length 3636
>>
stream
x�ŚkkG���W�Ǆ`4���`�c;6$�g7��A��:Y2����S5'�o��]���{W�u��\��l�sK�}�K��.M��ӻͶ����z[]Ҫw��x�EE=��������w�cIM�Җ4�nzO������1�R�e�1�'_~yr���������'��7�7o>?9����������{ϯ~>��鯯^]^�Ų�ܽ�]�~������'�nK���<{��p��m�NN���֓�Gg/^/M������W_vw�\�V<�!�Q�������������������[���A�1%:{yXN�y����_D{5����zqvm��\n����������E�+-��������ٽ�m������_�!��7�4:�������+���m�%�#W>�����޼��O.�v���Ã�[Yû������7���	+zga'�?-�u��U"�-��~)K]���]�FL)�5��K`T�+��z
�j��l{�(`џ1�WY�*$сw�Z�K��l� )��6�
����-Y߂�R�ء����/h@/R����4Mܳ���evA��,�O�Y�r�wո��"9L�c)�|M��5Ҩ�:�7靴�����S{�#��Wq"k�,�ʫ��Z��Ն8إA�ܒ`L��v��&vv�5��s�@�g^hk�{��6��j]
���Zu�H�º�V-Ucj{,[˚(4��C��3|s9h8m�ĸ��22���2���U\����M�ֹ�D�N؋
w��t-vݱVm�����}�������7V/�kJ���01qbךl�ԙ��F�_Lo�Ն�P��l�mS@�$6���B�^�S�"�EZ5ZIF��'�;8�ۀ!���0�:,�6�T*6��@��A!v��
� /I�I0�1�l��g���/��*���"[��_6h@y�⢽b�:WD��ތB�g�@I3hCCl�ȝ55�
�LL�:]%�!)�PG������%���kHY�hL`�)H�ٮv6-%-w��)�nJ��@)ŉN7	~VY�2�Z�r�@^qa�sU��.�pXy[�U%����L5^5�5���y�J�(/bH���}*�j���iȼ �FGֲf -t��;����֭L*U6���%���G��jG�w�n�Yp�lX��`P�"�W��%�ұ���9δ��K�0��L*��8߭
��;,A��Z����U�V�Z��fqu��o��nA��M�WO4 �Yg�;We���K	�/��%�a'�K�,�6���6x�/���f�bz���p��Zح��\숚z�ۑF���l�����bic���D_���Q=�z$�0���R�K�WF_��aTYXS��0��}������V��QQvL���X�!���5�5�h{��0�����sQ6؋��������Gr�)���\>E�p?�J�SEPD�h*��
%�Qx��m�+K��������:�G�u��2Ж�� �}3�6��?h���G✌�>��M ��dV>`[8�
�q{�w�m����B�w[p�חFðdZ`��x��C�41K3b��N�XE�j�B�	�S\�SM��m&�y?�@�̻�V����p���T=��(� ��HHn�ʛ$���WO�&��oT��>�"<
�4�¤&��*���x�_l�}Z�Tm[X2���J���L/��
�$�P�^5mu�:故��{\n��V������ش���*cT��&lP��ĉk��9M�Wa�k��O�Dv�::�"�ۻ��+FK5;���dTi8L;�n'\�Nw�&�vP��$����RXo�ܹ�.R��0�[/k�b��T*��a��³�̓J+ȯ1��c׈]�����H���(!JQQm���9���Aꞌ1<��F�ëJ5
�bYJ���Db�NBKvLu�Ȏ}�R�cFXM�1<� �۞�70�^��4��0b��{H9б�#���5y؛q��1k�-�߾�1+q�\��3X_D��߳C4�E��[.,�y�.!W�I݌=��]l��PG��N��4:���R�G�4$�!nL�lH#ƈ�� M�Tj��s5_�\���#��r8BL�2-#Ry˾U����f��OY�Y#����!��6�I��EO�Ֆ�i�D��h!�y�#��`6��L_7�V�IrD*�3�ٝ����U��:���X�H��y���.�u��Hx)Rg~"���օ�~x��[#pc�A������=��L�}�0ruYXP�X�S�D,MR�!<`��+��2E�]5�@G�":��K.�3|h�8��	�he����#?�{�j���h�!�Y�m�����@��}��<�0��m3�\��8y	���@vk$�>٫�m�6	��F�e�'�[�L?$�-I�L��M,�O���(1|*�X��`��f��C7卷V�Ev���%�Oω�+��u�BR��9Fns6x�t��f�wc*�40����3��8���;� jq�Y� ��H�%����&����AK��_bk�$?�� C���G!�H@���]cb޾�~��%D�rr'n䪄�n	;�"y�f��#F�n\���XgR����Dc`�d�\���L��ғ*�7W�Nú-�z�V��A�C�4kڤy�'��#�D+gG"57a�h�g��]?��)@?n+2jM���XFkn������[6�l;��F]
�!�
��"����7�d�p�����Y�|������2�Ԍ �zKҴ�i��3��g����NВp)Sǎ�7�UW|G�:N��R��Dp!�:X5��P$
�["��i��#qg��q����t�+�g?�ۓ�O�O ���8�1�3�
'!�0?.�����F�fu���8,p��Q���Y�n^Q���H�\�9�ɚǂ����q�2�p�8�3O���؇������3Ͻ~�>Y��E0������аq���U�#">��Aí!�V��Hǌ��CPu�:^��!;�Oq	��H�X�`�I���ƬeA^e�M�@�&Cٜ9�6?�-Z�Ṁ� ����Ѭ��qI�N�V߆� ��b���'f����7��GJ۩M��Ħm�8)��h�=7	������(����Z�^z�<�|v��۝���ΝǷn�WW�<WÃ�1�ݺT�bn]/�vw��w8��������섗h�����?a�����e���.���I�����?Nq�QKP��)���&$�������Ke<N���qA�%og��;�`��/G_�hW	8����5y��X���$��鏨���x���)rϠM�"��l0(N\��UA���8���T�q�%�����qɯ<N��lh��>~���/ه��}���e��Z
G��n,�o�޽�d���~��۳Wo��˶���i�s�9筋L�c�6��GrC�h~����>z�(̿�������n��7�)������f �����?�[�~�o!���<��Kp�w��{����?.����'�>��_����?���:��r��ՏW�"����1GL���3��o��Ͼ�w_.~y�𫯾{����ON�?���%mk<��h�
endstream
endobj
43 0 obj
<<
/Size 44
/Root 1 0 R
/Info 41 0 R
/ID [<05CEC68E3D92C0408099E91C2A165228> <74D8339AF50F2C0AF1E41FBFE5739311>]
/Type /XRef
/W [1 2 2]
/Filter /FlateDecode
/Index [0 44]
/Length 150
>>
stream
x�%�;
���]?�@�*^D;����,aA�Z����3X٬3$ŃdHֵU#��O�"x����PV}<0C�3�}��X$"���A&6�z�M�m��<��VW]��M�7�+�>%�))/�8��Y���/�?��
endstream
endobj
startxref
52095
%%EOF
